magic
tech sky130A
timestamp 1748436552
<< nwell >>
rect -87 331 160 491
<< pwell >>
rect -87 -19 160 100
<< scnmos >>
rect 60 24 75 89
<< scpmoshvt >>
rect 60 349 75 448
<< ndiff >>
rect 33 83 60 89
rect 33 66 37 83
rect 54 66 60 83
rect 33 49 60 66
rect 33 32 37 49
rect 54 32 60 49
rect 33 24 60 32
rect 75 83 102 89
rect 75 66 81 83
rect 98 66 102 83
rect 75 49 102 66
rect 75 32 81 49
rect 98 32 102 49
rect 75 24 102 32
<< pdiff >>
rect 33 442 60 448
rect 33 425 37 442
rect 54 425 60 442
rect 33 408 60 425
rect 33 391 37 408
rect 54 391 60 408
rect 33 374 60 391
rect 33 357 37 374
rect 54 357 60 374
rect 33 349 60 357
rect 75 442 102 448
rect 75 425 81 442
rect 98 425 102 442
rect 75 408 102 425
rect 75 391 81 408
rect 98 391 102 408
rect 75 374 102 391
rect 75 357 81 374
rect 98 357 102 374
rect 75 349 102 357
<< ndiffc >>
rect 37 66 54 83
rect 37 32 54 49
rect 81 66 98 83
rect 81 32 98 49
<< pdiffc >>
rect 37 425 54 442
rect 37 391 54 408
rect 37 357 54 374
rect 81 425 98 442
rect 81 391 98 408
rect 81 357 98 374
<< psubdiff >>
rect -34 77 6 89
rect -34 59 -20 77
rect -2 59 6 77
rect -34 24 6 59
<< nsubdiff >>
rect -34 379 6 448
rect -34 361 -16 379
rect 2 361 6 379
rect -34 349 6 361
<< psubdiffcont >>
rect -20 59 -2 77
<< nsubdiffcont >>
rect -16 361 2 379
<< poly >>
rect 60 448 75 461
rect 60 233 75 349
rect -87 226 75 233
rect -87 209 -75 226
rect -58 209 75 226
rect -87 201 75 209
rect 60 89 75 201
rect 60 11 75 24
<< polycont >>
rect -75 209 -58 226
<< locali >>
rect 0 463 14 481
rect 32 463 60 481
rect 78 463 106 481
rect 124 463 138 481
rect 31 442 54 463
rect 31 425 37 442
rect 31 408 54 425
rect 31 391 37 408
rect 31 387 54 391
rect -16 379 54 387
rect 2 374 54 379
rect 2 361 37 374
rect -16 357 37 361
rect -16 349 54 357
rect 72 442 106 446
rect 72 425 81 442
rect 98 425 106 442
rect 72 408 106 425
rect 72 391 81 408
rect 98 391 106 408
rect 72 374 106 391
rect 72 357 81 374
rect 98 357 106 374
rect 72 349 106 357
rect -87 226 -50 233
rect -87 209 -75 226
rect -58 209 -50 226
rect -87 201 -50 209
rect 81 228 106 349
rect 128 228 160 232
rect 81 227 160 228
rect 81 210 136 227
rect 153 210 160 227
rect 81 208 160 210
rect -33 83 54 91
rect 81 89 106 208
rect 128 204 160 208
rect -33 77 37 83
rect -33 59 -20 77
rect -2 66 37 77
rect -2 59 54 66
rect -33 55 54 59
rect 31 49 54 55
rect 31 32 37 49
rect 31 9 54 32
rect 72 83 106 89
rect 72 66 81 83
rect 98 66 106 83
rect 72 49 106 66
rect 72 32 81 49
rect 98 32 106 49
rect 72 26 106 32
rect 0 -9 14 9
rect 32 -9 60 9
rect 78 -9 106 9
rect 124 -9 138 9
<< viali >>
rect 14 463 32 481
rect 60 463 78 481
rect 106 463 124 481
rect -75 209 -58 226
rect 136 210 153 227
rect 14 -9 32 9
rect 60 -9 78 9
rect 106 -9 124 9
<< metal1 >>
rect -87 481 160 496
rect -87 463 14 481
rect 32 463 60 481
rect 78 463 106 481
rect 124 463 160 481
rect -87 448 160 463
rect -87 226 -50 233
rect -87 209 -75 226
rect -58 209 -50 226
rect -87 201 -50 209
rect 128 227 160 232
rect 128 210 136 227
rect 153 210 160 227
rect 128 204 160 210
rect -87 9 160 24
rect -87 -9 14 9
rect 32 -9 60 9
rect 78 -9 106 9
rect 124 -9 160 9
rect -87 -24 160 -9
<< labels >>
flabel metal1 -79 -12 -55 12 0 FreeSans 80 0 0 0 VGND
port 4 nsew power bidirectional
flabel metal1 -77 461 -53 485 0 FreeSans 80 0 0 0 VDPWR
port 5 nsew ground bidirectional
flabel metal1 -79 205 -55 229 0 FreeSans 80 0 0 0 A
port 8 nsew signal input
flabel metal1 133 206 157 230 0 FreeSans 80 0 0 0 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX -107 -44 180 316
string GDS_FILEBOUNDARY true
string LEFclass CORE
string LEForigin 0 0
string LEFsite unithd
<< end >>
