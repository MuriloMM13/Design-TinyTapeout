magic
tech sky130A
timestamp 1750757695
<< nwell >>
rect -87 331 160 592
<< pwell >>
rect -87 -23 160 100
<< scnmos >>
rect 60 24 75 89
<< scpmoshvt >>
rect 60 349 75 549
<< ndiff >>
rect 33 83 60 89
rect 33 66 37 83
rect 54 66 60 83
rect 33 49 60 66
rect 33 32 37 49
rect 54 32 60 49
rect 33 24 60 32
rect 75 83 102 89
rect 75 66 81 83
rect 98 66 102 83
rect 75 49 102 66
rect 75 32 81 49
rect 98 32 102 49
rect 75 24 102 32
<< pdiff >>
rect 33 526 60 549
rect 33 509 37 526
rect 54 509 60 526
rect 33 492 60 509
rect 33 475 37 492
rect 54 475 60 492
rect 33 458 60 475
rect 33 441 37 458
rect 54 441 60 458
rect 33 424 60 441
rect 33 407 37 424
rect 54 407 60 424
rect 33 390 60 407
rect 33 373 37 390
rect 54 373 60 390
rect 33 349 60 373
rect 75 526 102 549
rect 75 509 81 526
rect 98 509 102 526
rect 75 492 102 509
rect 75 475 81 492
rect 98 475 102 492
rect 75 458 102 475
rect 75 441 81 458
rect 98 441 102 458
rect 75 424 102 441
rect 75 407 81 424
rect 98 407 102 424
rect 75 390 102 407
rect 75 373 81 390
rect 98 373 102 390
rect 75 349 102 373
<< ndiffc >>
rect 37 66 54 83
rect 37 32 54 49
rect 81 66 98 83
rect 81 32 98 49
<< pdiffc >>
rect 37 509 54 526
rect 37 475 54 492
rect 37 441 54 458
rect 37 407 54 424
rect 37 373 54 390
rect 81 509 98 526
rect 81 475 98 492
rect 81 441 98 458
rect 81 407 98 424
rect 81 373 98 390
<< psubdiff >>
rect -34 77 6 89
rect -34 59 -20 77
rect -2 59 6 77
rect -34 24 6 59
<< nsubdiff >>
rect -34 379 6 549
rect -34 361 -16 379
rect 2 361 6 379
rect -34 349 6 361
<< psubdiffcont >>
rect -20 59 -2 77
<< nsubdiffcont >>
rect -16 361 2 379
<< poly >>
rect 60 549 75 562
rect -87 233 -39 241
rect 60 233 75 349
rect -87 226 75 233
rect -87 208 -72 226
rect -54 208 75 226
rect -87 201 75 208
rect -87 193 -39 201
rect 60 89 75 201
rect 60 11 75 24
<< polycont >>
rect -72 208 -54 226
<< locali >>
rect 0 564 14 582
rect 32 564 60 582
rect 78 564 106 582
rect 124 564 138 582
rect 31 526 54 564
rect 31 509 37 526
rect 31 492 54 509
rect 31 475 37 492
rect 31 458 54 475
rect 31 441 37 458
rect 31 424 54 441
rect 31 407 37 424
rect 31 390 54 407
rect 31 387 37 390
rect -16 379 37 387
rect 2 373 37 379
rect 2 361 54 373
rect -16 349 54 361
rect 72 526 106 534
rect 72 509 81 526
rect 98 509 106 526
rect 72 492 106 509
rect 72 475 81 492
rect 98 475 106 492
rect 72 458 106 475
rect 72 441 81 458
rect 98 441 106 458
rect 72 424 106 441
rect 72 407 81 424
rect 98 407 106 424
rect 72 390 106 407
rect 72 373 81 390
rect 98 373 106 390
rect 72 349 106 373
rect 81 242 106 349
rect -87 226 -39 241
rect -87 208 -72 226
rect -54 208 -39 226
rect -87 193 -39 208
rect 81 227 160 242
rect 81 209 121 227
rect 139 209 160 227
rect 81 194 160 209
rect -33 83 54 91
rect 81 89 106 194
rect -33 77 37 83
rect -33 59 -20 77
rect -2 66 37 77
rect -2 59 54 66
rect -33 55 54 59
rect 31 49 54 55
rect 31 32 37 49
rect 31 9 54 32
rect 72 83 106 89
rect 72 66 81 83
rect 98 66 106 83
rect 72 49 106 66
rect 72 32 81 49
rect 98 32 106 49
rect 72 26 106 32
rect 0 -9 14 9
rect 32 -9 60 9
rect 78 -9 106 9
rect 124 -9 138 9
<< viali >>
rect 14 564 32 582
rect 60 564 78 582
rect 106 564 124 582
rect -72 208 -54 226
rect 121 209 139 227
rect 14 -9 32 9
rect 60 -9 78 9
rect 106 -9 124 9
<< metal1 >>
rect -87 582 160 597
rect -87 564 14 582
rect 32 564 60 582
rect 78 564 106 582
rect 124 564 160 582
rect -87 549 160 564
rect -87 226 -39 241
rect -87 208 -72 226
rect -54 208 -39 226
rect -87 193 -39 208
rect 112 227 160 242
rect 112 209 121 227
rect 139 209 160 227
rect 112 194 160 209
rect -87 9 160 24
rect -87 -9 14 9
rect 32 -9 60 9
rect 78 -9 106 9
rect 124 -9 160 9
rect -87 -24 160 -9
<< labels >>
flabel metal1 -87 -24 -39 24 1 FreeSans 200 0 0 0 VGND
port 22 nsew ground bidirectional
flabel metal1 -87 193 -39 241 1 FreeSans 200 0 0 0 A
port 24 nsew signal input
flabel metal1 112 194 160 242 1 FreeSans 200 0 0 0 Y
port 25 nsew signal output
flabel metal1 -87 549 -39 597 1 FreeSans 200 0 0 0 VDPWR
port 23 nsew power bidirectional
<< properties >>
string FIXED_BBOX -107 -44 180 316
string GDS_FILEBOUNDARY true
string LEFclass CORE
string LEForigin 0 0
string LEFsite unithd
<< end >>
