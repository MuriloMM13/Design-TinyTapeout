VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mag/tt_um_analog_murilo
  CLASS BLOCK ;
  FOREIGN mag/tt_um_analog_murilo ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.010 BY 0.010 ;
END mag/tt_um_analog_murilo
END LIBRARY

