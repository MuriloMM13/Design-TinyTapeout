magic
tech sky130A
timestamp 1748162301
<< locali >>
rect 13259 971 13309 986
rect 15191 971 15241 986
rect 13259 970 14075 971
rect 13259 952 13275 970
rect 13293 952 14075 970
rect 13259 951 14075 952
rect 14254 970 15241 971
rect 14254 952 15207 970
rect 15225 952 15241 970
rect 14254 951 15241 952
rect 13259 936 13309 951
rect 15191 936 15241 951
<< viali >>
rect 13275 952 13293 970
rect 15207 952 15225 970
<< metal1 >>
rect 142 1139 192 1140
rect 142 1128 14075 1139
rect 142 1102 154 1128
rect 180 1102 14075 1128
rect 142 1091 14075 1102
rect 142 1090 192 1091
rect 13259 974 13309 986
rect 13259 948 13271 974
rect 13297 948 13309 974
rect 13259 936 13309 948
rect 15191 974 15241 986
rect 15191 948 15203 974
rect 15229 948 15241 974
rect 15191 936 15241 948
rect 448 867 498 868
rect 448 856 14075 867
rect 448 830 460 856
rect 486 830 14075 856
rect 448 819 14075 830
rect 448 818 498 819
<< via1 >>
rect 154 1102 180 1128
rect 13271 970 13297 974
rect 13271 952 13275 970
rect 13275 952 13293 970
rect 13293 952 13297 970
rect 13271 948 13297 952
rect 15203 970 15229 974
rect 15203 952 15207 970
rect 15207 952 15225 970
rect 15225 952 15229 970
rect 15203 948 15229 952
rect 460 830 486 856
<< metal2 >>
rect 142 1129 192 1140
rect 142 1101 153 1129
rect 181 1101 192 1129
rect 142 1090 192 1101
rect 13259 975 13309 986
rect 13259 947 13270 975
rect 13298 947 13309 975
rect 13259 936 13309 947
rect 15191 975 15241 986
rect 15191 947 15202 975
rect 15230 947 15241 975
rect 15191 936 15241 947
rect 448 857 498 868
rect 448 829 459 857
rect 487 829 498 857
rect 448 818 498 829
<< via2 >>
rect 153 1128 181 1129
rect 153 1102 154 1128
rect 154 1102 180 1128
rect 180 1102 181 1128
rect 153 1101 181 1102
rect 13270 974 13298 975
rect 13270 948 13271 974
rect 13271 948 13297 974
rect 13297 948 13298 974
rect 13270 947 13298 948
rect 15202 974 15230 975
rect 15202 948 15203 974
rect 15203 948 15229 974
rect 15229 948 15230 974
rect 15202 947 15230 948
rect 459 856 487 857
rect 459 830 460 856
rect 460 830 486 856
rect 486 830 487 856
rect 459 829 487 830
<< metal3 >>
rect 142 1131 192 1140
rect 142 1099 151 1131
rect 183 1099 192 1131
rect 142 1090 192 1099
rect 13259 977 13309 986
rect 13259 945 13268 977
rect 13300 945 13309 977
rect 13259 936 13309 945
rect 15191 977 15241 986
rect 15191 945 15200 977
rect 15232 945 15241 977
rect 15191 936 15241 945
rect 448 859 498 868
rect 448 827 457 859
rect 489 827 498 859
rect 448 818 498 827
<< via3 >>
rect 151 1129 183 1131
rect 151 1101 153 1129
rect 153 1101 181 1129
rect 181 1101 183 1129
rect 151 1099 183 1101
rect 13268 975 13300 977
rect 13268 947 13270 975
rect 13270 947 13298 975
rect 13298 947 13300 975
rect 13268 945 13300 947
rect 15200 975 15232 977
rect 15200 947 15202 975
rect 15202 947 15230 975
rect 15230 947 15232 975
rect 15200 945 15232 947
rect 457 857 489 859
rect 457 829 459 857
rect 459 829 487 857
rect 487 829 489 857
rect 457 827 489 829
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 7483 22476 7513 22576
rect 7759 22476 7789 22576
rect 8035 22476 8065 22576
rect 8311 22476 8341 22576
rect 8587 22476 8617 22576
rect 8863 22476 8893 22576
rect 9139 22476 9169 22576
rect 9415 22476 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 100 1131 300 22076
rect 100 1099 151 1131
rect 183 1099 300 1131
rect 100 500 300 1099
rect 400 859 600 22076
rect 400 827 457 859
rect 489 827 600 859
rect 400 500 600 827
rect 13249 977 13339 999
rect 13249 945 13268 977
rect 13300 945 13339 977
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 945
rect 15181 977 15271 999
rect 15181 945 15200 977
rect 15232 945 15271 977
rect 15181 0 15271 945
use NOT  NOT_0
timestamp 1748129733
transform 1 0 14094 0 1 843
box -81 -24 160 296
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 300 90 0 0 clk
port 1 nsew
flabel metal4 s 14398 22526 14398 22526 0 FreeSans 300 90 0 0 clk
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 300 90 0 0 ena
port 2 nsew
flabel metal4 s 14674 22526 14674 22526 0 FreeSans 300 90 0 0 ena
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 300 90 0 0 rst_n
port 3 nsew
flabel metal4 s 14122 22526 14122 22526 0 FreeSans 300 90 0 0 rst_n
flabel metal4 s 15181 0 15271 100 0 FreeSans 600 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 15226 50 15226 50 0 FreeSans 600 0 0 0 ua[0]
flabel metal4 s 13249 0 13339 100 0 FreeSans 600 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 13294 50 13294 50 0 FreeSans 600 0 0 0 ua[1]
flabel metal4 s 11317 0 11407 100 0 FreeSans 600 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 11362 50 11362 50 0 FreeSans 600 0 0 0 ua[2]
flabel metal4 s 9385 0 9475 100 0 FreeSans 600 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 9430 50 9430 50 0 FreeSans 600 0 0 0 ua[3]
flabel metal4 s 7453 0 7543 100 0 FreeSans 600 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 7498 50 7498 50 0 FreeSans 600 0 0 0 ua[4]
flabel metal4 s 5521 0 5611 100 0 FreeSans 600 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 5566 50 5566 50 0 FreeSans 600 0 0 0 ua[5]
flabel metal4 s 3589 0 3679 100 0 FreeSans 600 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 3634 50 3634 50 0 FreeSans 600 0 0 0 ua[6]
flabel metal4 s 1657 0 1747 100 0 FreeSans 600 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 1702 50 1702 50 0 FreeSans 600 0 0 0 ua[7]
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 300 90 0 0 ui_in[0]
port 12 nsew
flabel metal4 s 13846 22526 13846 22526 0 FreeSans 300 90 0 0 ui_in[0]
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 300 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 13570 22526 13570 22526 0 FreeSans 300 90 0 0 ui_in[1]
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 300 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 13294 22526 13294 22526 0 FreeSans 300 90 0 0 ui_in[2]
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 300 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 13018 22526 13018 22526 0 FreeSans 300 90 0 0 ui_in[3]
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 300 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 12742 22526 12742 22526 0 FreeSans 300 90 0 0 ui_in[4]
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 300 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 12466 22526 12466 22526 0 FreeSans 300 90 0 0 ui_in[5]
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 300 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 12190 22526 12190 22526 0 FreeSans 300 90 0 0 ui_in[6]
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 300 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 11914 22526 11914 22526 0 FreeSans 300 90 0 0 ui_in[7]
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 300 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 11638 22526 11638 22526 0 FreeSans 300 90 0 0 uio_in[0]
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 300 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 11362 22526 11362 22526 0 FreeSans 300 90 0 0 uio_in[1]
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 300 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 11086 22526 11086 22526 0 FreeSans 300 90 0 0 uio_in[2]
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 300 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 10810 22526 10810 22526 0 FreeSans 300 90 0 0 uio_in[3]
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 300 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 10534 22526 10534 22526 0 FreeSans 300 90 0 0 uio_in[4]
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 300 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 10258 22526 10258 22526 0 FreeSans 300 90 0 0 uio_in[5]
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 300 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 9982 22526 9982 22526 0 FreeSans 300 90 0 0 uio_in[6]
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 300 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 9706 22526 9706 22526 0 FreeSans 300 90 0 0 uio_in[7]
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 300 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 5014 22526 5014 22526 0 FreeSans 300 90 0 0 uio_oe[0]
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 300 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 4738 22526 4738 22526 0 FreeSans 300 90 0 0 uio_oe[1]
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 300 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 4462 22526 4462 22526 0 FreeSans 300 90 0 0 uio_oe[2]
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 300 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 4186 22526 4186 22526 0 FreeSans 300 90 0 0 uio_oe[3]
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 300 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 3910 22526 3910 22526 0 FreeSans 300 90 0 0 uio_oe[4]
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 300 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 3634 22526 3634 22526 0 FreeSans 300 90 0 0 uio_oe[5]
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 300 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 3358 22526 3358 22526 0 FreeSans 300 90 0 0 uio_oe[6]
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 300 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 3082 22526 3082 22526 0 FreeSans 300 90 0 0 uio_oe[7]
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 300 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 7222 22526 7222 22526 0 FreeSans 300 90 0 0 uio_out[0]
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 300 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 6946 22526 6946 22526 0 FreeSans 300 90 0 0 uio_out[1]
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 300 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 6670 22526 6670 22526 0 FreeSans 300 90 0 0 uio_out[2]
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 300 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 6394 22526 6394 22526 0 FreeSans 300 90 0 0 uio_out[3]
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 300 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 6118 22526 6118 22526 0 FreeSans 300 90 0 0 uio_out[4]
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 300 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 5842 22526 5842 22526 0 FreeSans 300 90 0 0 uio_out[5]
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 300 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 5566 22526 5566 22526 0 FreeSans 300 90 0 0 uio_out[6]
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 300 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 5290 22526 5290 22526 0 FreeSans 300 90 0 0 uio_out[7]
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 300 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 9430 22526 9430 22526 0 FreeSans 300 90 0 0 uo_out[0]
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 300 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 9154 22526 9154 22526 0 FreeSans 300 90 0 0 uo_out[1]
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 300 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 8878 22526 8878 22526 0 FreeSans 300 90 0 0 uo_out[2]
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 300 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 8602 22526 8602 22526 0 FreeSans 300 90 0 0 uo_out[3]
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 300 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 8326 22526 8326 22526 0 FreeSans 300 90 0 0 uo_out[4]
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 300 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 8050 22526 8050 22526 0 FreeSans 300 90 0 0 uo_out[5]
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 300 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 7774 22526 7774 22526 0 FreeSans 300 90 0 0 uo_out[6]
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 300 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 7498 22526 7498 22526 0 FreeSans 300 90 0 0 uo_out[7]
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 60 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 61 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
