VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOT
  CLASS CORE ;
  FOREIGN NOT ;
  ORIGIN 1.070 0.440 ;
  SIZE 2.870 BY 3.600 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.870 -0.240 -0.390 0.240 ;
    END
  END VGND
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.870 3.310 1.600 4.910 ;
      LAYER li1 ;
        RECT 0.000 4.630 1.380 4.810 ;
        RECT 0.310 3.870 0.540 4.630 ;
        RECT -0.160 3.490 0.540 3.870 ;
      LAYER met1 ;
        RECT -0.870 4.480 1.600 4.960 ;
    END
  END VDPWR
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER met1 ;
        RECT -0.870 1.930 -0.390 2.410 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.442800 ;
    PORT
      LAYER li1 ;
        RECT 0.720 3.490 1.060 4.460 ;
        RECT 0.810 3.160 1.060 3.490 ;
      LAYER met1 ;
        RECT 1.120 1.940 1.600 2.420 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT -0.870 -0.150 1.600 1.000 ;
        RECT -0.390 -0.190 1.600 -0.150 ;
      LAYER li1 ;
        RECT 0.810 2.420 1.060 3.160 ;
        RECT -0.870 1.930 -0.390 2.410 ;
        RECT 0.810 1.940 1.600 2.420 ;
        RECT -0.330 0.550 0.540 0.910 ;
        RECT 0.810 0.890 1.060 1.940 ;
        RECT 0.310 0.090 0.540 0.550 ;
        RECT 0.720 0.260 1.060 0.890 ;
        RECT 0.000 -0.090 1.380 0.090 ;
      LAYER met1 ;
        RECT -0.390 -0.240 1.600 0.240 ;
  END
END NOT
END LIBRARY

