magic
tech sky130A
timestamp 1753208556
<< nwell >>
rect 10113 7826 10286 8062
rect 10724 7826 10897 8062
rect 11302 7826 11475 8062
rect 11913 7826 12086 8062
rect 12524 7826 12697 8062
rect 9502 7176 9675 7412
rect 10113 7176 10286 7412
rect 10724 7176 10897 7412
rect 11302 7176 11475 7412
rect 11913 7176 12086 7412
rect 12524 7176 12697 7412
rect 9502 6536 9675 6772
rect 10113 6536 10286 6772
rect 10724 6536 10897 6772
rect 11302 6536 11475 6772
rect 11913 6536 12086 6772
rect 12524 6536 12697 6772
rect 9502 5886 9675 6122
rect 10113 5886 10286 6122
rect 10724 5886 10897 6122
rect 11302 5886 11475 6122
rect 11913 5886 12086 6122
rect 12524 5886 12697 6122
rect 9502 5236 9675 5472
rect 10113 5236 10286 5472
rect 10724 5236 10897 5472
rect 11302 5236 11475 5472
rect 11913 5236 12086 5472
rect 12524 5236 12697 5472
rect 9502 4596 9675 4832
rect 10113 4596 10286 4832
rect 10724 4596 10897 4832
rect 11302 4596 11475 4832
rect 11913 4596 12086 4832
rect 12524 4596 12697 4832
<< nmos >>
rect 10090 7570 10105 7670
rect 10126 7570 10141 7670
rect 10170 7570 10185 7670
rect 10214 7570 10229 7670
rect 10258 7570 10273 7670
rect 10294 7570 10309 7670
rect 10701 7570 10716 7670
rect 10737 7570 10752 7670
rect 10781 7570 10796 7670
rect 10825 7570 10840 7670
rect 10869 7570 10884 7670
rect 10905 7570 10920 7670
rect 11279 7570 11294 7670
rect 11315 7570 11330 7670
rect 11359 7570 11374 7670
rect 11403 7570 11418 7670
rect 11447 7570 11462 7670
rect 11483 7570 11498 7670
rect 11890 7570 11905 7670
rect 11926 7570 11941 7670
rect 11970 7570 11985 7670
rect 12014 7570 12029 7670
rect 12058 7570 12073 7670
rect 12094 7570 12109 7670
rect 12501 7570 12516 7670
rect 12537 7570 12552 7670
rect 12581 7570 12596 7670
rect 12625 7570 12640 7670
rect 12669 7570 12684 7670
rect 12705 7570 12720 7670
rect 9479 6920 9494 7020
rect 9515 6920 9530 7020
rect 9559 6920 9574 7020
rect 9603 6920 9618 7020
rect 9647 6920 9662 7020
rect 9683 6920 9698 7020
rect 10090 6920 10105 7020
rect 10126 6920 10141 7020
rect 10170 6920 10185 7020
rect 10214 6920 10229 7020
rect 10258 6920 10273 7020
rect 10294 6920 10309 7020
rect 10701 6920 10716 7020
rect 10737 6920 10752 7020
rect 10781 6920 10796 7020
rect 10825 6920 10840 7020
rect 10869 6920 10884 7020
rect 10905 6920 10920 7020
rect 11279 6920 11294 7020
rect 11315 6920 11330 7020
rect 11359 6920 11374 7020
rect 11403 6920 11418 7020
rect 11447 6920 11462 7020
rect 11483 6920 11498 7020
rect 11890 6920 11905 7020
rect 11926 6920 11941 7020
rect 11970 6920 11985 7020
rect 12014 6920 12029 7020
rect 12058 6920 12073 7020
rect 12094 6920 12109 7020
rect 12501 6920 12516 7020
rect 12537 6920 12552 7020
rect 12581 6920 12596 7020
rect 12625 6920 12640 7020
rect 12669 6920 12684 7020
rect 12705 6920 12720 7020
rect 9479 6280 9494 6380
rect 9515 6280 9530 6380
rect 9559 6280 9574 6380
rect 9603 6280 9618 6380
rect 9647 6280 9662 6380
rect 9683 6280 9698 6380
rect 10090 6280 10105 6380
rect 10126 6280 10141 6380
rect 10170 6280 10185 6380
rect 10214 6280 10229 6380
rect 10258 6280 10273 6380
rect 10294 6280 10309 6380
rect 10701 6280 10716 6380
rect 10737 6280 10752 6380
rect 10781 6280 10796 6380
rect 10825 6280 10840 6380
rect 10869 6280 10884 6380
rect 10905 6280 10920 6380
rect 11279 6280 11294 6380
rect 11315 6280 11330 6380
rect 11359 6280 11374 6380
rect 11403 6280 11418 6380
rect 11447 6280 11462 6380
rect 11483 6280 11498 6380
rect 11890 6280 11905 6380
rect 11926 6280 11941 6380
rect 11970 6280 11985 6380
rect 12014 6280 12029 6380
rect 12058 6280 12073 6380
rect 12094 6280 12109 6380
rect 12501 6280 12516 6380
rect 12537 6280 12552 6380
rect 12581 6280 12596 6380
rect 12625 6280 12640 6380
rect 12669 6280 12684 6380
rect 12705 6280 12720 6380
rect 9479 5630 9494 5730
rect 9515 5630 9530 5730
rect 9559 5630 9574 5730
rect 9603 5630 9618 5730
rect 9647 5630 9662 5730
rect 9683 5630 9698 5730
rect 10090 5630 10105 5730
rect 10126 5630 10141 5730
rect 10170 5630 10185 5730
rect 10214 5630 10229 5730
rect 10258 5630 10273 5730
rect 10294 5630 10309 5730
rect 10701 5630 10716 5730
rect 10737 5630 10752 5730
rect 10781 5630 10796 5730
rect 10825 5630 10840 5730
rect 10869 5630 10884 5730
rect 10905 5630 10920 5730
rect 11279 5630 11294 5730
rect 11315 5630 11330 5730
rect 11359 5630 11374 5730
rect 11403 5630 11418 5730
rect 11447 5630 11462 5730
rect 11483 5630 11498 5730
rect 11890 5630 11905 5730
rect 11926 5630 11941 5730
rect 11970 5630 11985 5730
rect 12014 5630 12029 5730
rect 12058 5630 12073 5730
rect 12094 5630 12109 5730
rect 12501 5630 12516 5730
rect 12537 5630 12552 5730
rect 12581 5630 12596 5730
rect 12625 5630 12640 5730
rect 12669 5630 12684 5730
rect 12705 5630 12720 5730
rect 9479 4980 9494 5080
rect 9515 4980 9530 5080
rect 9559 4980 9574 5080
rect 9603 4980 9618 5080
rect 9647 4980 9662 5080
rect 9683 4980 9698 5080
rect 10090 4980 10105 5080
rect 10126 4980 10141 5080
rect 10170 4980 10185 5080
rect 10214 4980 10229 5080
rect 10258 4980 10273 5080
rect 10294 4980 10309 5080
rect 10701 4980 10716 5080
rect 10737 4980 10752 5080
rect 10781 4980 10796 5080
rect 10825 4980 10840 5080
rect 10869 4980 10884 5080
rect 10905 4980 10920 5080
rect 11279 4980 11294 5080
rect 11315 4980 11330 5080
rect 11359 4980 11374 5080
rect 11403 4980 11418 5080
rect 11447 4980 11462 5080
rect 11483 4980 11498 5080
rect 11890 4980 11905 5080
rect 11926 4980 11941 5080
rect 11970 4980 11985 5080
rect 12014 4980 12029 5080
rect 12058 4980 12073 5080
rect 12094 4980 12109 5080
rect 12501 4980 12516 5080
rect 12537 4980 12552 5080
rect 12581 4980 12596 5080
rect 12625 4980 12640 5080
rect 12669 4980 12684 5080
rect 12705 4980 12720 5080
rect 9479 4340 9494 4440
rect 9515 4340 9530 4440
rect 9559 4340 9574 4440
rect 9603 4340 9618 4440
rect 9647 4340 9662 4440
rect 9683 4340 9698 4440
rect 10090 4340 10105 4440
rect 10126 4340 10141 4440
rect 10170 4340 10185 4440
rect 10214 4340 10229 4440
rect 10258 4340 10273 4440
rect 10294 4340 10309 4440
rect 10701 4340 10716 4440
rect 10737 4340 10752 4440
rect 10781 4340 10796 4440
rect 10825 4340 10840 4440
rect 10869 4340 10884 4440
rect 10905 4340 10920 4440
rect 11279 4340 11294 4440
rect 11315 4340 11330 4440
rect 11359 4340 11374 4440
rect 11403 4340 11418 4440
rect 11447 4340 11462 4440
rect 11483 4340 11498 4440
rect 11890 4340 11905 4440
rect 11926 4340 11941 4440
rect 11970 4340 11985 4440
rect 12014 4340 12029 4440
rect 12058 4340 12073 4440
rect 12094 4340 12109 4440
rect 12501 4340 12516 4440
rect 12537 4340 12552 4440
rect 12581 4340 12596 4440
rect 12625 4340 12640 4440
rect 12669 4340 12684 4440
rect 12705 4340 12720 4440
<< pmos >>
rect 10170 7844 10185 8044
rect 10214 7844 10229 8044
rect 10781 7844 10796 8044
rect 10825 7844 10840 8044
rect 11359 7844 11374 8044
rect 11403 7844 11418 8044
rect 11970 7844 11985 8044
rect 12014 7844 12029 8044
rect 12581 7844 12596 8044
rect 12625 7844 12640 8044
rect 9559 7194 9574 7394
rect 9603 7194 9618 7394
rect 10170 7194 10185 7394
rect 10214 7194 10229 7394
rect 10781 7194 10796 7394
rect 10825 7194 10840 7394
rect 11359 7194 11374 7394
rect 11403 7194 11418 7394
rect 11970 7194 11985 7394
rect 12014 7194 12029 7394
rect 12581 7194 12596 7394
rect 12625 7194 12640 7394
rect 9559 6554 9574 6754
rect 9603 6554 9618 6754
rect 10170 6554 10185 6754
rect 10214 6554 10229 6754
rect 10781 6554 10796 6754
rect 10825 6554 10840 6754
rect 11359 6554 11374 6754
rect 11403 6554 11418 6754
rect 11970 6554 11985 6754
rect 12014 6554 12029 6754
rect 12581 6554 12596 6754
rect 12625 6554 12640 6754
rect 9559 5904 9574 6104
rect 9603 5904 9618 6104
rect 10170 5904 10185 6104
rect 10214 5904 10229 6104
rect 10781 5904 10796 6104
rect 10825 5904 10840 6104
rect 11359 5904 11374 6104
rect 11403 5904 11418 6104
rect 11970 5904 11985 6104
rect 12014 5904 12029 6104
rect 12581 5904 12596 6104
rect 12625 5904 12640 6104
rect 9559 5254 9574 5454
rect 9603 5254 9618 5454
rect 10170 5254 10185 5454
rect 10214 5254 10229 5454
rect 10781 5254 10796 5454
rect 10825 5254 10840 5454
rect 11359 5254 11374 5454
rect 11403 5254 11418 5454
rect 11970 5254 11985 5454
rect 12014 5254 12029 5454
rect 12581 5254 12596 5454
rect 12625 5254 12640 5454
rect 9559 4614 9574 4814
rect 9603 4614 9618 4814
rect 10170 4614 10185 4814
rect 10214 4614 10229 4814
rect 10781 4614 10796 4814
rect 10825 4614 10840 4814
rect 11359 4614 11374 4814
rect 11403 4614 11418 4814
rect 11970 4614 11985 4814
rect 12014 4614 12029 4814
rect 12581 4614 12596 4814
rect 12625 4614 12640 4814
<< ndiff >>
rect 10061 7663 10090 7670
rect 10061 7646 10067 7663
rect 10084 7646 10090 7663
rect 10061 7629 10090 7646
rect 10061 7612 10067 7629
rect 10084 7612 10090 7629
rect 10061 7595 10090 7612
rect 10061 7578 10067 7595
rect 10084 7578 10090 7595
rect 10061 7570 10090 7578
rect 10105 7570 10126 7670
rect 10141 7663 10170 7670
rect 10141 7646 10147 7663
rect 10164 7646 10170 7663
rect 10141 7629 10170 7646
rect 10141 7612 10147 7629
rect 10164 7612 10170 7629
rect 10141 7595 10170 7612
rect 10141 7578 10147 7595
rect 10164 7578 10170 7595
rect 10141 7570 10170 7578
rect 10185 7663 10214 7670
rect 10185 7646 10191 7663
rect 10208 7646 10214 7663
rect 10185 7629 10214 7646
rect 10185 7612 10191 7629
rect 10208 7612 10214 7629
rect 10185 7595 10214 7612
rect 10185 7578 10191 7595
rect 10208 7578 10214 7595
rect 10185 7570 10214 7578
rect 10229 7663 10258 7670
rect 10229 7646 10235 7663
rect 10252 7646 10258 7663
rect 10229 7629 10258 7646
rect 10229 7612 10235 7629
rect 10252 7612 10258 7629
rect 10229 7595 10258 7612
rect 10229 7578 10235 7595
rect 10252 7578 10258 7595
rect 10229 7570 10258 7578
rect 10273 7570 10294 7670
rect 10309 7663 10338 7670
rect 10309 7646 10315 7663
rect 10332 7646 10338 7663
rect 10309 7629 10338 7646
rect 10309 7612 10315 7629
rect 10332 7612 10338 7629
rect 10309 7595 10338 7612
rect 10309 7578 10315 7595
rect 10332 7578 10338 7595
rect 10309 7570 10338 7578
rect 10672 7663 10701 7670
rect 10672 7646 10678 7663
rect 10695 7646 10701 7663
rect 10672 7629 10701 7646
rect 10672 7612 10678 7629
rect 10695 7612 10701 7629
rect 10672 7595 10701 7612
rect 10672 7578 10678 7595
rect 10695 7578 10701 7595
rect 10672 7570 10701 7578
rect 10716 7570 10737 7670
rect 10752 7663 10781 7670
rect 10752 7646 10758 7663
rect 10775 7646 10781 7663
rect 10752 7629 10781 7646
rect 10752 7612 10758 7629
rect 10775 7612 10781 7629
rect 10752 7595 10781 7612
rect 10752 7578 10758 7595
rect 10775 7578 10781 7595
rect 10752 7570 10781 7578
rect 10796 7663 10825 7670
rect 10796 7646 10802 7663
rect 10819 7646 10825 7663
rect 10796 7629 10825 7646
rect 10796 7612 10802 7629
rect 10819 7612 10825 7629
rect 10796 7595 10825 7612
rect 10796 7578 10802 7595
rect 10819 7578 10825 7595
rect 10796 7570 10825 7578
rect 10840 7663 10869 7670
rect 10840 7646 10846 7663
rect 10863 7646 10869 7663
rect 10840 7629 10869 7646
rect 10840 7612 10846 7629
rect 10863 7612 10869 7629
rect 10840 7595 10869 7612
rect 10840 7578 10846 7595
rect 10863 7578 10869 7595
rect 10840 7570 10869 7578
rect 10884 7570 10905 7670
rect 10920 7663 10949 7670
rect 10920 7646 10926 7663
rect 10943 7646 10949 7663
rect 10920 7629 10949 7646
rect 10920 7612 10926 7629
rect 10943 7612 10949 7629
rect 10920 7595 10949 7612
rect 10920 7578 10926 7595
rect 10943 7578 10949 7595
rect 10920 7570 10949 7578
rect 11250 7663 11279 7670
rect 11250 7646 11256 7663
rect 11273 7646 11279 7663
rect 11250 7629 11279 7646
rect 11250 7612 11256 7629
rect 11273 7612 11279 7629
rect 11250 7595 11279 7612
rect 11250 7578 11256 7595
rect 11273 7578 11279 7595
rect 11250 7570 11279 7578
rect 11294 7570 11315 7670
rect 11330 7663 11359 7670
rect 11330 7646 11336 7663
rect 11353 7646 11359 7663
rect 11330 7629 11359 7646
rect 11330 7612 11336 7629
rect 11353 7612 11359 7629
rect 11330 7595 11359 7612
rect 11330 7578 11336 7595
rect 11353 7578 11359 7595
rect 11330 7570 11359 7578
rect 11374 7663 11403 7670
rect 11374 7646 11380 7663
rect 11397 7646 11403 7663
rect 11374 7629 11403 7646
rect 11374 7612 11380 7629
rect 11397 7612 11403 7629
rect 11374 7595 11403 7612
rect 11374 7578 11380 7595
rect 11397 7578 11403 7595
rect 11374 7570 11403 7578
rect 11418 7663 11447 7670
rect 11418 7646 11424 7663
rect 11441 7646 11447 7663
rect 11418 7629 11447 7646
rect 11418 7612 11424 7629
rect 11441 7612 11447 7629
rect 11418 7595 11447 7612
rect 11418 7578 11424 7595
rect 11441 7578 11447 7595
rect 11418 7570 11447 7578
rect 11462 7570 11483 7670
rect 11498 7663 11527 7670
rect 11498 7646 11504 7663
rect 11521 7646 11527 7663
rect 11498 7629 11527 7646
rect 11498 7612 11504 7629
rect 11521 7612 11527 7629
rect 11498 7595 11527 7612
rect 11498 7578 11504 7595
rect 11521 7578 11527 7595
rect 11498 7570 11527 7578
rect 11861 7663 11890 7670
rect 11861 7646 11867 7663
rect 11884 7646 11890 7663
rect 11861 7629 11890 7646
rect 11861 7612 11867 7629
rect 11884 7612 11890 7629
rect 11861 7595 11890 7612
rect 11861 7578 11867 7595
rect 11884 7578 11890 7595
rect 11861 7570 11890 7578
rect 11905 7570 11926 7670
rect 11941 7663 11970 7670
rect 11941 7646 11947 7663
rect 11964 7646 11970 7663
rect 11941 7629 11970 7646
rect 11941 7612 11947 7629
rect 11964 7612 11970 7629
rect 11941 7595 11970 7612
rect 11941 7578 11947 7595
rect 11964 7578 11970 7595
rect 11941 7570 11970 7578
rect 11985 7663 12014 7670
rect 11985 7646 11991 7663
rect 12008 7646 12014 7663
rect 11985 7629 12014 7646
rect 11985 7612 11991 7629
rect 12008 7612 12014 7629
rect 11985 7595 12014 7612
rect 11985 7578 11991 7595
rect 12008 7578 12014 7595
rect 11985 7570 12014 7578
rect 12029 7663 12058 7670
rect 12029 7646 12035 7663
rect 12052 7646 12058 7663
rect 12029 7629 12058 7646
rect 12029 7612 12035 7629
rect 12052 7612 12058 7629
rect 12029 7595 12058 7612
rect 12029 7578 12035 7595
rect 12052 7578 12058 7595
rect 12029 7570 12058 7578
rect 12073 7570 12094 7670
rect 12109 7663 12138 7670
rect 12109 7646 12115 7663
rect 12132 7646 12138 7663
rect 12109 7629 12138 7646
rect 12109 7612 12115 7629
rect 12132 7612 12138 7629
rect 12109 7595 12138 7612
rect 12109 7578 12115 7595
rect 12132 7578 12138 7595
rect 12109 7570 12138 7578
rect 12472 7663 12501 7670
rect 12472 7646 12478 7663
rect 12495 7646 12501 7663
rect 12472 7629 12501 7646
rect 12472 7612 12478 7629
rect 12495 7612 12501 7629
rect 12472 7595 12501 7612
rect 12472 7578 12478 7595
rect 12495 7578 12501 7595
rect 12472 7570 12501 7578
rect 12516 7570 12537 7670
rect 12552 7663 12581 7670
rect 12552 7646 12558 7663
rect 12575 7646 12581 7663
rect 12552 7629 12581 7646
rect 12552 7612 12558 7629
rect 12575 7612 12581 7629
rect 12552 7595 12581 7612
rect 12552 7578 12558 7595
rect 12575 7578 12581 7595
rect 12552 7570 12581 7578
rect 12596 7663 12625 7670
rect 12596 7646 12602 7663
rect 12619 7646 12625 7663
rect 12596 7629 12625 7646
rect 12596 7612 12602 7629
rect 12619 7612 12625 7629
rect 12596 7595 12625 7612
rect 12596 7578 12602 7595
rect 12619 7578 12625 7595
rect 12596 7570 12625 7578
rect 12640 7663 12669 7670
rect 12640 7646 12646 7663
rect 12663 7646 12669 7663
rect 12640 7629 12669 7646
rect 12640 7612 12646 7629
rect 12663 7612 12669 7629
rect 12640 7595 12669 7612
rect 12640 7578 12646 7595
rect 12663 7578 12669 7595
rect 12640 7570 12669 7578
rect 12684 7570 12705 7670
rect 12720 7663 12749 7670
rect 12720 7646 12726 7663
rect 12743 7646 12749 7663
rect 12720 7629 12749 7646
rect 12720 7612 12726 7629
rect 12743 7612 12749 7629
rect 12720 7595 12749 7612
rect 12720 7578 12726 7595
rect 12743 7578 12749 7595
rect 12720 7570 12749 7578
rect 9450 7013 9479 7020
rect 9450 6996 9456 7013
rect 9473 6996 9479 7013
rect 9450 6979 9479 6996
rect 9450 6962 9456 6979
rect 9473 6962 9479 6979
rect 9450 6945 9479 6962
rect 9450 6928 9456 6945
rect 9473 6928 9479 6945
rect 9450 6920 9479 6928
rect 9494 6920 9515 7020
rect 9530 7013 9559 7020
rect 9530 6996 9536 7013
rect 9553 6996 9559 7013
rect 9530 6979 9559 6996
rect 9530 6962 9536 6979
rect 9553 6962 9559 6979
rect 9530 6945 9559 6962
rect 9530 6928 9536 6945
rect 9553 6928 9559 6945
rect 9530 6920 9559 6928
rect 9574 7013 9603 7020
rect 9574 6996 9580 7013
rect 9597 6996 9603 7013
rect 9574 6979 9603 6996
rect 9574 6962 9580 6979
rect 9597 6962 9603 6979
rect 9574 6945 9603 6962
rect 9574 6928 9580 6945
rect 9597 6928 9603 6945
rect 9574 6920 9603 6928
rect 9618 7013 9647 7020
rect 9618 6996 9624 7013
rect 9641 6996 9647 7013
rect 9618 6979 9647 6996
rect 9618 6962 9624 6979
rect 9641 6962 9647 6979
rect 9618 6945 9647 6962
rect 9618 6928 9624 6945
rect 9641 6928 9647 6945
rect 9618 6920 9647 6928
rect 9662 6920 9683 7020
rect 9698 7013 9727 7020
rect 9698 6996 9704 7013
rect 9721 6996 9727 7013
rect 9698 6979 9727 6996
rect 9698 6962 9704 6979
rect 9721 6962 9727 6979
rect 9698 6945 9727 6962
rect 9698 6928 9704 6945
rect 9721 6928 9727 6945
rect 9698 6920 9727 6928
rect 10061 7013 10090 7020
rect 10061 6996 10067 7013
rect 10084 6996 10090 7013
rect 10061 6979 10090 6996
rect 10061 6962 10067 6979
rect 10084 6962 10090 6979
rect 10061 6945 10090 6962
rect 10061 6928 10067 6945
rect 10084 6928 10090 6945
rect 10061 6920 10090 6928
rect 10105 6920 10126 7020
rect 10141 7013 10170 7020
rect 10141 6996 10147 7013
rect 10164 6996 10170 7013
rect 10141 6979 10170 6996
rect 10141 6962 10147 6979
rect 10164 6962 10170 6979
rect 10141 6945 10170 6962
rect 10141 6928 10147 6945
rect 10164 6928 10170 6945
rect 10141 6920 10170 6928
rect 10185 7013 10214 7020
rect 10185 6996 10191 7013
rect 10208 6996 10214 7013
rect 10185 6979 10214 6996
rect 10185 6962 10191 6979
rect 10208 6962 10214 6979
rect 10185 6945 10214 6962
rect 10185 6928 10191 6945
rect 10208 6928 10214 6945
rect 10185 6920 10214 6928
rect 10229 7013 10258 7020
rect 10229 6996 10235 7013
rect 10252 6996 10258 7013
rect 10229 6979 10258 6996
rect 10229 6962 10235 6979
rect 10252 6962 10258 6979
rect 10229 6945 10258 6962
rect 10229 6928 10235 6945
rect 10252 6928 10258 6945
rect 10229 6920 10258 6928
rect 10273 6920 10294 7020
rect 10309 7013 10338 7020
rect 10309 6996 10315 7013
rect 10332 6996 10338 7013
rect 10309 6979 10338 6996
rect 10309 6962 10315 6979
rect 10332 6962 10338 6979
rect 10309 6945 10338 6962
rect 10309 6928 10315 6945
rect 10332 6928 10338 6945
rect 10309 6920 10338 6928
rect 10672 7013 10701 7020
rect 10672 6996 10678 7013
rect 10695 6996 10701 7013
rect 10672 6979 10701 6996
rect 10672 6962 10678 6979
rect 10695 6962 10701 6979
rect 10672 6945 10701 6962
rect 10672 6928 10678 6945
rect 10695 6928 10701 6945
rect 10672 6920 10701 6928
rect 10716 6920 10737 7020
rect 10752 7013 10781 7020
rect 10752 6996 10758 7013
rect 10775 6996 10781 7013
rect 10752 6979 10781 6996
rect 10752 6962 10758 6979
rect 10775 6962 10781 6979
rect 10752 6945 10781 6962
rect 10752 6928 10758 6945
rect 10775 6928 10781 6945
rect 10752 6920 10781 6928
rect 10796 7013 10825 7020
rect 10796 6996 10802 7013
rect 10819 6996 10825 7013
rect 10796 6979 10825 6996
rect 10796 6962 10802 6979
rect 10819 6962 10825 6979
rect 10796 6945 10825 6962
rect 10796 6928 10802 6945
rect 10819 6928 10825 6945
rect 10796 6920 10825 6928
rect 10840 7013 10869 7020
rect 10840 6996 10846 7013
rect 10863 6996 10869 7013
rect 10840 6979 10869 6996
rect 10840 6962 10846 6979
rect 10863 6962 10869 6979
rect 10840 6945 10869 6962
rect 10840 6928 10846 6945
rect 10863 6928 10869 6945
rect 10840 6920 10869 6928
rect 10884 6920 10905 7020
rect 10920 7013 10949 7020
rect 10920 6996 10926 7013
rect 10943 6996 10949 7013
rect 10920 6979 10949 6996
rect 10920 6962 10926 6979
rect 10943 6962 10949 6979
rect 10920 6945 10949 6962
rect 10920 6928 10926 6945
rect 10943 6928 10949 6945
rect 10920 6920 10949 6928
rect 11250 7013 11279 7020
rect 11250 6996 11256 7013
rect 11273 6996 11279 7013
rect 11250 6979 11279 6996
rect 11250 6962 11256 6979
rect 11273 6962 11279 6979
rect 11250 6945 11279 6962
rect 11250 6928 11256 6945
rect 11273 6928 11279 6945
rect 11250 6920 11279 6928
rect 11294 6920 11315 7020
rect 11330 7013 11359 7020
rect 11330 6996 11336 7013
rect 11353 6996 11359 7013
rect 11330 6979 11359 6996
rect 11330 6962 11336 6979
rect 11353 6962 11359 6979
rect 11330 6945 11359 6962
rect 11330 6928 11336 6945
rect 11353 6928 11359 6945
rect 11330 6920 11359 6928
rect 11374 7013 11403 7020
rect 11374 6996 11380 7013
rect 11397 6996 11403 7013
rect 11374 6979 11403 6996
rect 11374 6962 11380 6979
rect 11397 6962 11403 6979
rect 11374 6945 11403 6962
rect 11374 6928 11380 6945
rect 11397 6928 11403 6945
rect 11374 6920 11403 6928
rect 11418 7013 11447 7020
rect 11418 6996 11424 7013
rect 11441 6996 11447 7013
rect 11418 6979 11447 6996
rect 11418 6962 11424 6979
rect 11441 6962 11447 6979
rect 11418 6945 11447 6962
rect 11418 6928 11424 6945
rect 11441 6928 11447 6945
rect 11418 6920 11447 6928
rect 11462 6920 11483 7020
rect 11498 7013 11527 7020
rect 11498 6996 11504 7013
rect 11521 6996 11527 7013
rect 11498 6979 11527 6996
rect 11498 6962 11504 6979
rect 11521 6962 11527 6979
rect 11498 6945 11527 6962
rect 11498 6928 11504 6945
rect 11521 6928 11527 6945
rect 11498 6920 11527 6928
rect 11861 7013 11890 7020
rect 11861 6996 11867 7013
rect 11884 6996 11890 7013
rect 11861 6979 11890 6996
rect 11861 6962 11867 6979
rect 11884 6962 11890 6979
rect 11861 6945 11890 6962
rect 11861 6928 11867 6945
rect 11884 6928 11890 6945
rect 11861 6920 11890 6928
rect 11905 6920 11926 7020
rect 11941 7013 11970 7020
rect 11941 6996 11947 7013
rect 11964 6996 11970 7013
rect 11941 6979 11970 6996
rect 11941 6962 11947 6979
rect 11964 6962 11970 6979
rect 11941 6945 11970 6962
rect 11941 6928 11947 6945
rect 11964 6928 11970 6945
rect 11941 6920 11970 6928
rect 11985 7013 12014 7020
rect 11985 6996 11991 7013
rect 12008 6996 12014 7013
rect 11985 6979 12014 6996
rect 11985 6962 11991 6979
rect 12008 6962 12014 6979
rect 11985 6945 12014 6962
rect 11985 6928 11991 6945
rect 12008 6928 12014 6945
rect 11985 6920 12014 6928
rect 12029 7013 12058 7020
rect 12029 6996 12035 7013
rect 12052 6996 12058 7013
rect 12029 6979 12058 6996
rect 12029 6962 12035 6979
rect 12052 6962 12058 6979
rect 12029 6945 12058 6962
rect 12029 6928 12035 6945
rect 12052 6928 12058 6945
rect 12029 6920 12058 6928
rect 12073 6920 12094 7020
rect 12109 7013 12138 7020
rect 12109 6996 12115 7013
rect 12132 6996 12138 7013
rect 12109 6979 12138 6996
rect 12109 6962 12115 6979
rect 12132 6962 12138 6979
rect 12109 6945 12138 6962
rect 12109 6928 12115 6945
rect 12132 6928 12138 6945
rect 12109 6920 12138 6928
rect 12472 7013 12501 7020
rect 12472 6996 12478 7013
rect 12495 6996 12501 7013
rect 12472 6979 12501 6996
rect 12472 6962 12478 6979
rect 12495 6962 12501 6979
rect 12472 6945 12501 6962
rect 12472 6928 12478 6945
rect 12495 6928 12501 6945
rect 12472 6920 12501 6928
rect 12516 6920 12537 7020
rect 12552 7013 12581 7020
rect 12552 6996 12558 7013
rect 12575 6996 12581 7013
rect 12552 6979 12581 6996
rect 12552 6962 12558 6979
rect 12575 6962 12581 6979
rect 12552 6945 12581 6962
rect 12552 6928 12558 6945
rect 12575 6928 12581 6945
rect 12552 6920 12581 6928
rect 12596 7013 12625 7020
rect 12596 6996 12602 7013
rect 12619 6996 12625 7013
rect 12596 6979 12625 6996
rect 12596 6962 12602 6979
rect 12619 6962 12625 6979
rect 12596 6945 12625 6962
rect 12596 6928 12602 6945
rect 12619 6928 12625 6945
rect 12596 6920 12625 6928
rect 12640 7013 12669 7020
rect 12640 6996 12646 7013
rect 12663 6996 12669 7013
rect 12640 6979 12669 6996
rect 12640 6962 12646 6979
rect 12663 6962 12669 6979
rect 12640 6945 12669 6962
rect 12640 6928 12646 6945
rect 12663 6928 12669 6945
rect 12640 6920 12669 6928
rect 12684 6920 12705 7020
rect 12720 7013 12749 7020
rect 12720 6996 12726 7013
rect 12743 6996 12749 7013
rect 12720 6979 12749 6996
rect 12720 6962 12726 6979
rect 12743 6962 12749 6979
rect 12720 6945 12749 6962
rect 12720 6928 12726 6945
rect 12743 6928 12749 6945
rect 12720 6920 12749 6928
rect 9450 6373 9479 6380
rect 9450 6356 9456 6373
rect 9473 6356 9479 6373
rect 9450 6339 9479 6356
rect 9450 6322 9456 6339
rect 9473 6322 9479 6339
rect 9450 6305 9479 6322
rect 9450 6288 9456 6305
rect 9473 6288 9479 6305
rect 9450 6280 9479 6288
rect 9494 6280 9515 6380
rect 9530 6373 9559 6380
rect 9530 6356 9536 6373
rect 9553 6356 9559 6373
rect 9530 6339 9559 6356
rect 9530 6322 9536 6339
rect 9553 6322 9559 6339
rect 9530 6305 9559 6322
rect 9530 6288 9536 6305
rect 9553 6288 9559 6305
rect 9530 6280 9559 6288
rect 9574 6373 9603 6380
rect 9574 6356 9580 6373
rect 9597 6356 9603 6373
rect 9574 6339 9603 6356
rect 9574 6322 9580 6339
rect 9597 6322 9603 6339
rect 9574 6305 9603 6322
rect 9574 6288 9580 6305
rect 9597 6288 9603 6305
rect 9574 6280 9603 6288
rect 9618 6373 9647 6380
rect 9618 6356 9624 6373
rect 9641 6356 9647 6373
rect 9618 6339 9647 6356
rect 9618 6322 9624 6339
rect 9641 6322 9647 6339
rect 9618 6305 9647 6322
rect 9618 6288 9624 6305
rect 9641 6288 9647 6305
rect 9618 6280 9647 6288
rect 9662 6280 9683 6380
rect 9698 6373 9727 6380
rect 9698 6356 9704 6373
rect 9721 6356 9727 6373
rect 9698 6339 9727 6356
rect 9698 6322 9704 6339
rect 9721 6322 9727 6339
rect 9698 6305 9727 6322
rect 9698 6288 9704 6305
rect 9721 6288 9727 6305
rect 9698 6280 9727 6288
rect 10061 6373 10090 6380
rect 10061 6356 10067 6373
rect 10084 6356 10090 6373
rect 10061 6339 10090 6356
rect 10061 6322 10067 6339
rect 10084 6322 10090 6339
rect 10061 6305 10090 6322
rect 10061 6288 10067 6305
rect 10084 6288 10090 6305
rect 10061 6280 10090 6288
rect 10105 6280 10126 6380
rect 10141 6373 10170 6380
rect 10141 6356 10147 6373
rect 10164 6356 10170 6373
rect 10141 6339 10170 6356
rect 10141 6322 10147 6339
rect 10164 6322 10170 6339
rect 10141 6305 10170 6322
rect 10141 6288 10147 6305
rect 10164 6288 10170 6305
rect 10141 6280 10170 6288
rect 10185 6373 10214 6380
rect 10185 6356 10191 6373
rect 10208 6356 10214 6373
rect 10185 6339 10214 6356
rect 10185 6322 10191 6339
rect 10208 6322 10214 6339
rect 10185 6305 10214 6322
rect 10185 6288 10191 6305
rect 10208 6288 10214 6305
rect 10185 6280 10214 6288
rect 10229 6373 10258 6380
rect 10229 6356 10235 6373
rect 10252 6356 10258 6373
rect 10229 6339 10258 6356
rect 10229 6322 10235 6339
rect 10252 6322 10258 6339
rect 10229 6305 10258 6322
rect 10229 6288 10235 6305
rect 10252 6288 10258 6305
rect 10229 6280 10258 6288
rect 10273 6280 10294 6380
rect 10309 6373 10338 6380
rect 10309 6356 10315 6373
rect 10332 6356 10338 6373
rect 10309 6339 10338 6356
rect 10309 6322 10315 6339
rect 10332 6322 10338 6339
rect 10309 6305 10338 6322
rect 10309 6288 10315 6305
rect 10332 6288 10338 6305
rect 10309 6280 10338 6288
rect 10672 6373 10701 6380
rect 10672 6356 10678 6373
rect 10695 6356 10701 6373
rect 10672 6339 10701 6356
rect 10672 6322 10678 6339
rect 10695 6322 10701 6339
rect 10672 6305 10701 6322
rect 10672 6288 10678 6305
rect 10695 6288 10701 6305
rect 10672 6280 10701 6288
rect 10716 6280 10737 6380
rect 10752 6373 10781 6380
rect 10752 6356 10758 6373
rect 10775 6356 10781 6373
rect 10752 6339 10781 6356
rect 10752 6322 10758 6339
rect 10775 6322 10781 6339
rect 10752 6305 10781 6322
rect 10752 6288 10758 6305
rect 10775 6288 10781 6305
rect 10752 6280 10781 6288
rect 10796 6373 10825 6380
rect 10796 6356 10802 6373
rect 10819 6356 10825 6373
rect 10796 6339 10825 6356
rect 10796 6322 10802 6339
rect 10819 6322 10825 6339
rect 10796 6305 10825 6322
rect 10796 6288 10802 6305
rect 10819 6288 10825 6305
rect 10796 6280 10825 6288
rect 10840 6373 10869 6380
rect 10840 6356 10846 6373
rect 10863 6356 10869 6373
rect 10840 6339 10869 6356
rect 10840 6322 10846 6339
rect 10863 6322 10869 6339
rect 10840 6305 10869 6322
rect 10840 6288 10846 6305
rect 10863 6288 10869 6305
rect 10840 6280 10869 6288
rect 10884 6280 10905 6380
rect 10920 6373 10949 6380
rect 10920 6356 10926 6373
rect 10943 6356 10949 6373
rect 10920 6339 10949 6356
rect 10920 6322 10926 6339
rect 10943 6322 10949 6339
rect 10920 6305 10949 6322
rect 10920 6288 10926 6305
rect 10943 6288 10949 6305
rect 10920 6280 10949 6288
rect 11250 6373 11279 6380
rect 11250 6356 11256 6373
rect 11273 6356 11279 6373
rect 11250 6339 11279 6356
rect 11250 6322 11256 6339
rect 11273 6322 11279 6339
rect 11250 6305 11279 6322
rect 11250 6288 11256 6305
rect 11273 6288 11279 6305
rect 11250 6280 11279 6288
rect 11294 6280 11315 6380
rect 11330 6373 11359 6380
rect 11330 6356 11336 6373
rect 11353 6356 11359 6373
rect 11330 6339 11359 6356
rect 11330 6322 11336 6339
rect 11353 6322 11359 6339
rect 11330 6305 11359 6322
rect 11330 6288 11336 6305
rect 11353 6288 11359 6305
rect 11330 6280 11359 6288
rect 11374 6373 11403 6380
rect 11374 6356 11380 6373
rect 11397 6356 11403 6373
rect 11374 6339 11403 6356
rect 11374 6322 11380 6339
rect 11397 6322 11403 6339
rect 11374 6305 11403 6322
rect 11374 6288 11380 6305
rect 11397 6288 11403 6305
rect 11374 6280 11403 6288
rect 11418 6373 11447 6380
rect 11418 6356 11424 6373
rect 11441 6356 11447 6373
rect 11418 6339 11447 6356
rect 11418 6322 11424 6339
rect 11441 6322 11447 6339
rect 11418 6305 11447 6322
rect 11418 6288 11424 6305
rect 11441 6288 11447 6305
rect 11418 6280 11447 6288
rect 11462 6280 11483 6380
rect 11498 6373 11527 6380
rect 11498 6356 11504 6373
rect 11521 6356 11527 6373
rect 11498 6339 11527 6356
rect 11498 6322 11504 6339
rect 11521 6322 11527 6339
rect 11498 6305 11527 6322
rect 11498 6288 11504 6305
rect 11521 6288 11527 6305
rect 11498 6280 11527 6288
rect 11861 6373 11890 6380
rect 11861 6356 11867 6373
rect 11884 6356 11890 6373
rect 11861 6339 11890 6356
rect 11861 6322 11867 6339
rect 11884 6322 11890 6339
rect 11861 6305 11890 6322
rect 11861 6288 11867 6305
rect 11884 6288 11890 6305
rect 11861 6280 11890 6288
rect 11905 6280 11926 6380
rect 11941 6373 11970 6380
rect 11941 6356 11947 6373
rect 11964 6356 11970 6373
rect 11941 6339 11970 6356
rect 11941 6322 11947 6339
rect 11964 6322 11970 6339
rect 11941 6305 11970 6322
rect 11941 6288 11947 6305
rect 11964 6288 11970 6305
rect 11941 6280 11970 6288
rect 11985 6373 12014 6380
rect 11985 6356 11991 6373
rect 12008 6356 12014 6373
rect 11985 6339 12014 6356
rect 11985 6322 11991 6339
rect 12008 6322 12014 6339
rect 11985 6305 12014 6322
rect 11985 6288 11991 6305
rect 12008 6288 12014 6305
rect 11985 6280 12014 6288
rect 12029 6373 12058 6380
rect 12029 6356 12035 6373
rect 12052 6356 12058 6373
rect 12029 6339 12058 6356
rect 12029 6322 12035 6339
rect 12052 6322 12058 6339
rect 12029 6305 12058 6322
rect 12029 6288 12035 6305
rect 12052 6288 12058 6305
rect 12029 6280 12058 6288
rect 12073 6280 12094 6380
rect 12109 6373 12138 6380
rect 12109 6356 12115 6373
rect 12132 6356 12138 6373
rect 12109 6339 12138 6356
rect 12109 6322 12115 6339
rect 12132 6322 12138 6339
rect 12109 6305 12138 6322
rect 12109 6288 12115 6305
rect 12132 6288 12138 6305
rect 12109 6280 12138 6288
rect 12472 6373 12501 6380
rect 12472 6356 12478 6373
rect 12495 6356 12501 6373
rect 12472 6339 12501 6356
rect 12472 6322 12478 6339
rect 12495 6322 12501 6339
rect 12472 6305 12501 6322
rect 12472 6288 12478 6305
rect 12495 6288 12501 6305
rect 12472 6280 12501 6288
rect 12516 6280 12537 6380
rect 12552 6373 12581 6380
rect 12552 6356 12558 6373
rect 12575 6356 12581 6373
rect 12552 6339 12581 6356
rect 12552 6322 12558 6339
rect 12575 6322 12581 6339
rect 12552 6305 12581 6322
rect 12552 6288 12558 6305
rect 12575 6288 12581 6305
rect 12552 6280 12581 6288
rect 12596 6373 12625 6380
rect 12596 6356 12602 6373
rect 12619 6356 12625 6373
rect 12596 6339 12625 6356
rect 12596 6322 12602 6339
rect 12619 6322 12625 6339
rect 12596 6305 12625 6322
rect 12596 6288 12602 6305
rect 12619 6288 12625 6305
rect 12596 6280 12625 6288
rect 12640 6373 12669 6380
rect 12640 6356 12646 6373
rect 12663 6356 12669 6373
rect 12640 6339 12669 6356
rect 12640 6322 12646 6339
rect 12663 6322 12669 6339
rect 12640 6305 12669 6322
rect 12640 6288 12646 6305
rect 12663 6288 12669 6305
rect 12640 6280 12669 6288
rect 12684 6280 12705 6380
rect 12720 6373 12749 6380
rect 12720 6356 12726 6373
rect 12743 6356 12749 6373
rect 12720 6339 12749 6356
rect 12720 6322 12726 6339
rect 12743 6322 12749 6339
rect 12720 6305 12749 6322
rect 12720 6288 12726 6305
rect 12743 6288 12749 6305
rect 12720 6280 12749 6288
rect 9450 5723 9479 5730
rect 9450 5706 9456 5723
rect 9473 5706 9479 5723
rect 9450 5689 9479 5706
rect 9450 5672 9456 5689
rect 9473 5672 9479 5689
rect 9450 5655 9479 5672
rect 9450 5638 9456 5655
rect 9473 5638 9479 5655
rect 9450 5630 9479 5638
rect 9494 5630 9515 5730
rect 9530 5723 9559 5730
rect 9530 5706 9536 5723
rect 9553 5706 9559 5723
rect 9530 5689 9559 5706
rect 9530 5672 9536 5689
rect 9553 5672 9559 5689
rect 9530 5655 9559 5672
rect 9530 5638 9536 5655
rect 9553 5638 9559 5655
rect 9530 5630 9559 5638
rect 9574 5723 9603 5730
rect 9574 5706 9580 5723
rect 9597 5706 9603 5723
rect 9574 5689 9603 5706
rect 9574 5672 9580 5689
rect 9597 5672 9603 5689
rect 9574 5655 9603 5672
rect 9574 5638 9580 5655
rect 9597 5638 9603 5655
rect 9574 5630 9603 5638
rect 9618 5723 9647 5730
rect 9618 5706 9624 5723
rect 9641 5706 9647 5723
rect 9618 5689 9647 5706
rect 9618 5672 9624 5689
rect 9641 5672 9647 5689
rect 9618 5655 9647 5672
rect 9618 5638 9624 5655
rect 9641 5638 9647 5655
rect 9618 5630 9647 5638
rect 9662 5630 9683 5730
rect 9698 5723 9727 5730
rect 9698 5706 9704 5723
rect 9721 5706 9727 5723
rect 9698 5689 9727 5706
rect 9698 5672 9704 5689
rect 9721 5672 9727 5689
rect 9698 5655 9727 5672
rect 9698 5638 9704 5655
rect 9721 5638 9727 5655
rect 9698 5630 9727 5638
rect 10061 5723 10090 5730
rect 10061 5706 10067 5723
rect 10084 5706 10090 5723
rect 10061 5689 10090 5706
rect 10061 5672 10067 5689
rect 10084 5672 10090 5689
rect 10061 5655 10090 5672
rect 10061 5638 10067 5655
rect 10084 5638 10090 5655
rect 10061 5630 10090 5638
rect 10105 5630 10126 5730
rect 10141 5723 10170 5730
rect 10141 5706 10147 5723
rect 10164 5706 10170 5723
rect 10141 5689 10170 5706
rect 10141 5672 10147 5689
rect 10164 5672 10170 5689
rect 10141 5655 10170 5672
rect 10141 5638 10147 5655
rect 10164 5638 10170 5655
rect 10141 5630 10170 5638
rect 10185 5723 10214 5730
rect 10185 5706 10191 5723
rect 10208 5706 10214 5723
rect 10185 5689 10214 5706
rect 10185 5672 10191 5689
rect 10208 5672 10214 5689
rect 10185 5655 10214 5672
rect 10185 5638 10191 5655
rect 10208 5638 10214 5655
rect 10185 5630 10214 5638
rect 10229 5723 10258 5730
rect 10229 5706 10235 5723
rect 10252 5706 10258 5723
rect 10229 5689 10258 5706
rect 10229 5672 10235 5689
rect 10252 5672 10258 5689
rect 10229 5655 10258 5672
rect 10229 5638 10235 5655
rect 10252 5638 10258 5655
rect 10229 5630 10258 5638
rect 10273 5630 10294 5730
rect 10309 5723 10338 5730
rect 10309 5706 10315 5723
rect 10332 5706 10338 5723
rect 10309 5689 10338 5706
rect 10309 5672 10315 5689
rect 10332 5672 10338 5689
rect 10309 5655 10338 5672
rect 10309 5638 10315 5655
rect 10332 5638 10338 5655
rect 10309 5630 10338 5638
rect 10672 5723 10701 5730
rect 10672 5706 10678 5723
rect 10695 5706 10701 5723
rect 10672 5689 10701 5706
rect 10672 5672 10678 5689
rect 10695 5672 10701 5689
rect 10672 5655 10701 5672
rect 10672 5638 10678 5655
rect 10695 5638 10701 5655
rect 10672 5630 10701 5638
rect 10716 5630 10737 5730
rect 10752 5723 10781 5730
rect 10752 5706 10758 5723
rect 10775 5706 10781 5723
rect 10752 5689 10781 5706
rect 10752 5672 10758 5689
rect 10775 5672 10781 5689
rect 10752 5655 10781 5672
rect 10752 5638 10758 5655
rect 10775 5638 10781 5655
rect 10752 5630 10781 5638
rect 10796 5723 10825 5730
rect 10796 5706 10802 5723
rect 10819 5706 10825 5723
rect 10796 5689 10825 5706
rect 10796 5672 10802 5689
rect 10819 5672 10825 5689
rect 10796 5655 10825 5672
rect 10796 5638 10802 5655
rect 10819 5638 10825 5655
rect 10796 5630 10825 5638
rect 10840 5723 10869 5730
rect 10840 5706 10846 5723
rect 10863 5706 10869 5723
rect 10840 5689 10869 5706
rect 10840 5672 10846 5689
rect 10863 5672 10869 5689
rect 10840 5655 10869 5672
rect 10840 5638 10846 5655
rect 10863 5638 10869 5655
rect 10840 5630 10869 5638
rect 10884 5630 10905 5730
rect 10920 5723 10949 5730
rect 10920 5706 10926 5723
rect 10943 5706 10949 5723
rect 10920 5689 10949 5706
rect 10920 5672 10926 5689
rect 10943 5672 10949 5689
rect 10920 5655 10949 5672
rect 10920 5638 10926 5655
rect 10943 5638 10949 5655
rect 10920 5630 10949 5638
rect 11250 5723 11279 5730
rect 11250 5706 11256 5723
rect 11273 5706 11279 5723
rect 11250 5689 11279 5706
rect 11250 5672 11256 5689
rect 11273 5672 11279 5689
rect 11250 5655 11279 5672
rect 11250 5638 11256 5655
rect 11273 5638 11279 5655
rect 11250 5630 11279 5638
rect 11294 5630 11315 5730
rect 11330 5723 11359 5730
rect 11330 5706 11336 5723
rect 11353 5706 11359 5723
rect 11330 5689 11359 5706
rect 11330 5672 11336 5689
rect 11353 5672 11359 5689
rect 11330 5655 11359 5672
rect 11330 5638 11336 5655
rect 11353 5638 11359 5655
rect 11330 5630 11359 5638
rect 11374 5723 11403 5730
rect 11374 5706 11380 5723
rect 11397 5706 11403 5723
rect 11374 5689 11403 5706
rect 11374 5672 11380 5689
rect 11397 5672 11403 5689
rect 11374 5655 11403 5672
rect 11374 5638 11380 5655
rect 11397 5638 11403 5655
rect 11374 5630 11403 5638
rect 11418 5723 11447 5730
rect 11418 5706 11424 5723
rect 11441 5706 11447 5723
rect 11418 5689 11447 5706
rect 11418 5672 11424 5689
rect 11441 5672 11447 5689
rect 11418 5655 11447 5672
rect 11418 5638 11424 5655
rect 11441 5638 11447 5655
rect 11418 5630 11447 5638
rect 11462 5630 11483 5730
rect 11498 5723 11527 5730
rect 11498 5706 11504 5723
rect 11521 5706 11527 5723
rect 11498 5689 11527 5706
rect 11498 5672 11504 5689
rect 11521 5672 11527 5689
rect 11498 5655 11527 5672
rect 11498 5638 11504 5655
rect 11521 5638 11527 5655
rect 11498 5630 11527 5638
rect 11861 5723 11890 5730
rect 11861 5706 11867 5723
rect 11884 5706 11890 5723
rect 11861 5689 11890 5706
rect 11861 5672 11867 5689
rect 11884 5672 11890 5689
rect 11861 5655 11890 5672
rect 11861 5638 11867 5655
rect 11884 5638 11890 5655
rect 11861 5630 11890 5638
rect 11905 5630 11926 5730
rect 11941 5723 11970 5730
rect 11941 5706 11947 5723
rect 11964 5706 11970 5723
rect 11941 5689 11970 5706
rect 11941 5672 11947 5689
rect 11964 5672 11970 5689
rect 11941 5655 11970 5672
rect 11941 5638 11947 5655
rect 11964 5638 11970 5655
rect 11941 5630 11970 5638
rect 11985 5723 12014 5730
rect 11985 5706 11991 5723
rect 12008 5706 12014 5723
rect 11985 5689 12014 5706
rect 11985 5672 11991 5689
rect 12008 5672 12014 5689
rect 11985 5655 12014 5672
rect 11985 5638 11991 5655
rect 12008 5638 12014 5655
rect 11985 5630 12014 5638
rect 12029 5723 12058 5730
rect 12029 5706 12035 5723
rect 12052 5706 12058 5723
rect 12029 5689 12058 5706
rect 12029 5672 12035 5689
rect 12052 5672 12058 5689
rect 12029 5655 12058 5672
rect 12029 5638 12035 5655
rect 12052 5638 12058 5655
rect 12029 5630 12058 5638
rect 12073 5630 12094 5730
rect 12109 5723 12138 5730
rect 12109 5706 12115 5723
rect 12132 5706 12138 5723
rect 12109 5689 12138 5706
rect 12109 5672 12115 5689
rect 12132 5672 12138 5689
rect 12109 5655 12138 5672
rect 12109 5638 12115 5655
rect 12132 5638 12138 5655
rect 12109 5630 12138 5638
rect 12472 5723 12501 5730
rect 12472 5706 12478 5723
rect 12495 5706 12501 5723
rect 12472 5689 12501 5706
rect 12472 5672 12478 5689
rect 12495 5672 12501 5689
rect 12472 5655 12501 5672
rect 12472 5638 12478 5655
rect 12495 5638 12501 5655
rect 12472 5630 12501 5638
rect 12516 5630 12537 5730
rect 12552 5723 12581 5730
rect 12552 5706 12558 5723
rect 12575 5706 12581 5723
rect 12552 5689 12581 5706
rect 12552 5672 12558 5689
rect 12575 5672 12581 5689
rect 12552 5655 12581 5672
rect 12552 5638 12558 5655
rect 12575 5638 12581 5655
rect 12552 5630 12581 5638
rect 12596 5723 12625 5730
rect 12596 5706 12602 5723
rect 12619 5706 12625 5723
rect 12596 5689 12625 5706
rect 12596 5672 12602 5689
rect 12619 5672 12625 5689
rect 12596 5655 12625 5672
rect 12596 5638 12602 5655
rect 12619 5638 12625 5655
rect 12596 5630 12625 5638
rect 12640 5723 12669 5730
rect 12640 5706 12646 5723
rect 12663 5706 12669 5723
rect 12640 5689 12669 5706
rect 12640 5672 12646 5689
rect 12663 5672 12669 5689
rect 12640 5655 12669 5672
rect 12640 5638 12646 5655
rect 12663 5638 12669 5655
rect 12640 5630 12669 5638
rect 12684 5630 12705 5730
rect 12720 5723 12749 5730
rect 12720 5706 12726 5723
rect 12743 5706 12749 5723
rect 12720 5689 12749 5706
rect 12720 5672 12726 5689
rect 12743 5672 12749 5689
rect 12720 5655 12749 5672
rect 12720 5638 12726 5655
rect 12743 5638 12749 5655
rect 12720 5630 12749 5638
rect 9450 5073 9479 5080
rect 9450 5056 9456 5073
rect 9473 5056 9479 5073
rect 9450 5039 9479 5056
rect 9450 5022 9456 5039
rect 9473 5022 9479 5039
rect 9450 5005 9479 5022
rect 9450 4988 9456 5005
rect 9473 4988 9479 5005
rect 9450 4980 9479 4988
rect 9494 4980 9515 5080
rect 9530 5073 9559 5080
rect 9530 5056 9536 5073
rect 9553 5056 9559 5073
rect 9530 5039 9559 5056
rect 9530 5022 9536 5039
rect 9553 5022 9559 5039
rect 9530 5005 9559 5022
rect 9530 4988 9536 5005
rect 9553 4988 9559 5005
rect 9530 4980 9559 4988
rect 9574 5073 9603 5080
rect 9574 5056 9580 5073
rect 9597 5056 9603 5073
rect 9574 5039 9603 5056
rect 9574 5022 9580 5039
rect 9597 5022 9603 5039
rect 9574 5005 9603 5022
rect 9574 4988 9580 5005
rect 9597 4988 9603 5005
rect 9574 4980 9603 4988
rect 9618 5073 9647 5080
rect 9618 5056 9624 5073
rect 9641 5056 9647 5073
rect 9618 5039 9647 5056
rect 9618 5022 9624 5039
rect 9641 5022 9647 5039
rect 9618 5005 9647 5022
rect 9618 4988 9624 5005
rect 9641 4988 9647 5005
rect 9618 4980 9647 4988
rect 9662 4980 9683 5080
rect 9698 5073 9727 5080
rect 9698 5056 9704 5073
rect 9721 5056 9727 5073
rect 9698 5039 9727 5056
rect 9698 5022 9704 5039
rect 9721 5022 9727 5039
rect 9698 5005 9727 5022
rect 9698 4988 9704 5005
rect 9721 4988 9727 5005
rect 9698 4980 9727 4988
rect 10061 5073 10090 5080
rect 10061 5056 10067 5073
rect 10084 5056 10090 5073
rect 10061 5039 10090 5056
rect 10061 5022 10067 5039
rect 10084 5022 10090 5039
rect 10061 5005 10090 5022
rect 10061 4988 10067 5005
rect 10084 4988 10090 5005
rect 10061 4980 10090 4988
rect 10105 4980 10126 5080
rect 10141 5073 10170 5080
rect 10141 5056 10147 5073
rect 10164 5056 10170 5073
rect 10141 5039 10170 5056
rect 10141 5022 10147 5039
rect 10164 5022 10170 5039
rect 10141 5005 10170 5022
rect 10141 4988 10147 5005
rect 10164 4988 10170 5005
rect 10141 4980 10170 4988
rect 10185 5073 10214 5080
rect 10185 5056 10191 5073
rect 10208 5056 10214 5073
rect 10185 5039 10214 5056
rect 10185 5022 10191 5039
rect 10208 5022 10214 5039
rect 10185 5005 10214 5022
rect 10185 4988 10191 5005
rect 10208 4988 10214 5005
rect 10185 4980 10214 4988
rect 10229 5073 10258 5080
rect 10229 5056 10235 5073
rect 10252 5056 10258 5073
rect 10229 5039 10258 5056
rect 10229 5022 10235 5039
rect 10252 5022 10258 5039
rect 10229 5005 10258 5022
rect 10229 4988 10235 5005
rect 10252 4988 10258 5005
rect 10229 4980 10258 4988
rect 10273 4980 10294 5080
rect 10309 5073 10338 5080
rect 10309 5056 10315 5073
rect 10332 5056 10338 5073
rect 10309 5039 10338 5056
rect 10309 5022 10315 5039
rect 10332 5022 10338 5039
rect 10309 5005 10338 5022
rect 10309 4988 10315 5005
rect 10332 4988 10338 5005
rect 10309 4980 10338 4988
rect 10672 5073 10701 5080
rect 10672 5056 10678 5073
rect 10695 5056 10701 5073
rect 10672 5039 10701 5056
rect 10672 5022 10678 5039
rect 10695 5022 10701 5039
rect 10672 5005 10701 5022
rect 10672 4988 10678 5005
rect 10695 4988 10701 5005
rect 10672 4980 10701 4988
rect 10716 4980 10737 5080
rect 10752 5073 10781 5080
rect 10752 5056 10758 5073
rect 10775 5056 10781 5073
rect 10752 5039 10781 5056
rect 10752 5022 10758 5039
rect 10775 5022 10781 5039
rect 10752 5005 10781 5022
rect 10752 4988 10758 5005
rect 10775 4988 10781 5005
rect 10752 4980 10781 4988
rect 10796 5073 10825 5080
rect 10796 5056 10802 5073
rect 10819 5056 10825 5073
rect 10796 5039 10825 5056
rect 10796 5022 10802 5039
rect 10819 5022 10825 5039
rect 10796 5005 10825 5022
rect 10796 4988 10802 5005
rect 10819 4988 10825 5005
rect 10796 4980 10825 4988
rect 10840 5073 10869 5080
rect 10840 5056 10846 5073
rect 10863 5056 10869 5073
rect 10840 5039 10869 5056
rect 10840 5022 10846 5039
rect 10863 5022 10869 5039
rect 10840 5005 10869 5022
rect 10840 4988 10846 5005
rect 10863 4988 10869 5005
rect 10840 4980 10869 4988
rect 10884 4980 10905 5080
rect 10920 5073 10949 5080
rect 10920 5056 10926 5073
rect 10943 5056 10949 5073
rect 10920 5039 10949 5056
rect 10920 5022 10926 5039
rect 10943 5022 10949 5039
rect 10920 5005 10949 5022
rect 10920 4988 10926 5005
rect 10943 4988 10949 5005
rect 10920 4980 10949 4988
rect 11250 5073 11279 5080
rect 11250 5056 11256 5073
rect 11273 5056 11279 5073
rect 11250 5039 11279 5056
rect 11250 5022 11256 5039
rect 11273 5022 11279 5039
rect 11250 5005 11279 5022
rect 11250 4988 11256 5005
rect 11273 4988 11279 5005
rect 11250 4980 11279 4988
rect 11294 4980 11315 5080
rect 11330 5073 11359 5080
rect 11330 5056 11336 5073
rect 11353 5056 11359 5073
rect 11330 5039 11359 5056
rect 11330 5022 11336 5039
rect 11353 5022 11359 5039
rect 11330 5005 11359 5022
rect 11330 4988 11336 5005
rect 11353 4988 11359 5005
rect 11330 4980 11359 4988
rect 11374 5073 11403 5080
rect 11374 5056 11380 5073
rect 11397 5056 11403 5073
rect 11374 5039 11403 5056
rect 11374 5022 11380 5039
rect 11397 5022 11403 5039
rect 11374 5005 11403 5022
rect 11374 4988 11380 5005
rect 11397 4988 11403 5005
rect 11374 4980 11403 4988
rect 11418 5073 11447 5080
rect 11418 5056 11424 5073
rect 11441 5056 11447 5073
rect 11418 5039 11447 5056
rect 11418 5022 11424 5039
rect 11441 5022 11447 5039
rect 11418 5005 11447 5022
rect 11418 4988 11424 5005
rect 11441 4988 11447 5005
rect 11418 4980 11447 4988
rect 11462 4980 11483 5080
rect 11498 5073 11527 5080
rect 11498 5056 11504 5073
rect 11521 5056 11527 5073
rect 11498 5039 11527 5056
rect 11498 5022 11504 5039
rect 11521 5022 11527 5039
rect 11498 5005 11527 5022
rect 11498 4988 11504 5005
rect 11521 4988 11527 5005
rect 11498 4980 11527 4988
rect 11861 5073 11890 5080
rect 11861 5056 11867 5073
rect 11884 5056 11890 5073
rect 11861 5039 11890 5056
rect 11861 5022 11867 5039
rect 11884 5022 11890 5039
rect 11861 5005 11890 5022
rect 11861 4988 11867 5005
rect 11884 4988 11890 5005
rect 11861 4980 11890 4988
rect 11905 4980 11926 5080
rect 11941 5073 11970 5080
rect 11941 5056 11947 5073
rect 11964 5056 11970 5073
rect 11941 5039 11970 5056
rect 11941 5022 11947 5039
rect 11964 5022 11970 5039
rect 11941 5005 11970 5022
rect 11941 4988 11947 5005
rect 11964 4988 11970 5005
rect 11941 4980 11970 4988
rect 11985 5073 12014 5080
rect 11985 5056 11991 5073
rect 12008 5056 12014 5073
rect 11985 5039 12014 5056
rect 11985 5022 11991 5039
rect 12008 5022 12014 5039
rect 11985 5005 12014 5022
rect 11985 4988 11991 5005
rect 12008 4988 12014 5005
rect 11985 4980 12014 4988
rect 12029 5073 12058 5080
rect 12029 5056 12035 5073
rect 12052 5056 12058 5073
rect 12029 5039 12058 5056
rect 12029 5022 12035 5039
rect 12052 5022 12058 5039
rect 12029 5005 12058 5022
rect 12029 4988 12035 5005
rect 12052 4988 12058 5005
rect 12029 4980 12058 4988
rect 12073 4980 12094 5080
rect 12109 5073 12138 5080
rect 12109 5056 12115 5073
rect 12132 5056 12138 5073
rect 12109 5039 12138 5056
rect 12109 5022 12115 5039
rect 12132 5022 12138 5039
rect 12109 5005 12138 5022
rect 12109 4988 12115 5005
rect 12132 4988 12138 5005
rect 12109 4980 12138 4988
rect 12472 5073 12501 5080
rect 12472 5056 12478 5073
rect 12495 5056 12501 5073
rect 12472 5039 12501 5056
rect 12472 5022 12478 5039
rect 12495 5022 12501 5039
rect 12472 5005 12501 5022
rect 12472 4988 12478 5005
rect 12495 4988 12501 5005
rect 12472 4980 12501 4988
rect 12516 4980 12537 5080
rect 12552 5073 12581 5080
rect 12552 5056 12558 5073
rect 12575 5056 12581 5073
rect 12552 5039 12581 5056
rect 12552 5022 12558 5039
rect 12575 5022 12581 5039
rect 12552 5005 12581 5022
rect 12552 4988 12558 5005
rect 12575 4988 12581 5005
rect 12552 4980 12581 4988
rect 12596 5073 12625 5080
rect 12596 5056 12602 5073
rect 12619 5056 12625 5073
rect 12596 5039 12625 5056
rect 12596 5022 12602 5039
rect 12619 5022 12625 5039
rect 12596 5005 12625 5022
rect 12596 4988 12602 5005
rect 12619 4988 12625 5005
rect 12596 4980 12625 4988
rect 12640 5073 12669 5080
rect 12640 5056 12646 5073
rect 12663 5056 12669 5073
rect 12640 5039 12669 5056
rect 12640 5022 12646 5039
rect 12663 5022 12669 5039
rect 12640 5005 12669 5022
rect 12640 4988 12646 5005
rect 12663 4988 12669 5005
rect 12640 4980 12669 4988
rect 12684 4980 12705 5080
rect 12720 5073 12749 5080
rect 12720 5056 12726 5073
rect 12743 5056 12749 5073
rect 12720 5039 12749 5056
rect 12720 5022 12726 5039
rect 12743 5022 12749 5039
rect 12720 5005 12749 5022
rect 12720 4988 12726 5005
rect 12743 4988 12749 5005
rect 12720 4980 12749 4988
rect 9450 4433 9479 4440
rect 9450 4416 9456 4433
rect 9473 4416 9479 4433
rect 9450 4399 9479 4416
rect 9450 4382 9456 4399
rect 9473 4382 9479 4399
rect 9450 4365 9479 4382
rect 9450 4348 9456 4365
rect 9473 4348 9479 4365
rect 9450 4340 9479 4348
rect 9494 4340 9515 4440
rect 9530 4433 9559 4440
rect 9530 4416 9536 4433
rect 9553 4416 9559 4433
rect 9530 4399 9559 4416
rect 9530 4382 9536 4399
rect 9553 4382 9559 4399
rect 9530 4365 9559 4382
rect 9530 4348 9536 4365
rect 9553 4348 9559 4365
rect 9530 4340 9559 4348
rect 9574 4433 9603 4440
rect 9574 4416 9580 4433
rect 9597 4416 9603 4433
rect 9574 4399 9603 4416
rect 9574 4382 9580 4399
rect 9597 4382 9603 4399
rect 9574 4365 9603 4382
rect 9574 4348 9580 4365
rect 9597 4348 9603 4365
rect 9574 4340 9603 4348
rect 9618 4433 9647 4440
rect 9618 4416 9624 4433
rect 9641 4416 9647 4433
rect 9618 4399 9647 4416
rect 9618 4382 9624 4399
rect 9641 4382 9647 4399
rect 9618 4365 9647 4382
rect 9618 4348 9624 4365
rect 9641 4348 9647 4365
rect 9618 4340 9647 4348
rect 9662 4340 9683 4440
rect 9698 4433 9727 4440
rect 9698 4416 9704 4433
rect 9721 4416 9727 4433
rect 9698 4399 9727 4416
rect 9698 4382 9704 4399
rect 9721 4382 9727 4399
rect 9698 4365 9727 4382
rect 9698 4348 9704 4365
rect 9721 4348 9727 4365
rect 9698 4340 9727 4348
rect 10061 4433 10090 4440
rect 10061 4416 10067 4433
rect 10084 4416 10090 4433
rect 10061 4399 10090 4416
rect 10061 4382 10067 4399
rect 10084 4382 10090 4399
rect 10061 4365 10090 4382
rect 10061 4348 10067 4365
rect 10084 4348 10090 4365
rect 10061 4340 10090 4348
rect 10105 4340 10126 4440
rect 10141 4433 10170 4440
rect 10141 4416 10147 4433
rect 10164 4416 10170 4433
rect 10141 4399 10170 4416
rect 10141 4382 10147 4399
rect 10164 4382 10170 4399
rect 10141 4365 10170 4382
rect 10141 4348 10147 4365
rect 10164 4348 10170 4365
rect 10141 4340 10170 4348
rect 10185 4433 10214 4440
rect 10185 4416 10191 4433
rect 10208 4416 10214 4433
rect 10185 4399 10214 4416
rect 10185 4382 10191 4399
rect 10208 4382 10214 4399
rect 10185 4365 10214 4382
rect 10185 4348 10191 4365
rect 10208 4348 10214 4365
rect 10185 4340 10214 4348
rect 10229 4433 10258 4440
rect 10229 4416 10235 4433
rect 10252 4416 10258 4433
rect 10229 4399 10258 4416
rect 10229 4382 10235 4399
rect 10252 4382 10258 4399
rect 10229 4365 10258 4382
rect 10229 4348 10235 4365
rect 10252 4348 10258 4365
rect 10229 4340 10258 4348
rect 10273 4340 10294 4440
rect 10309 4433 10338 4440
rect 10309 4416 10315 4433
rect 10332 4416 10338 4433
rect 10309 4399 10338 4416
rect 10309 4382 10315 4399
rect 10332 4382 10338 4399
rect 10309 4365 10338 4382
rect 10309 4348 10315 4365
rect 10332 4348 10338 4365
rect 10309 4340 10338 4348
rect 10672 4433 10701 4440
rect 10672 4416 10678 4433
rect 10695 4416 10701 4433
rect 10672 4399 10701 4416
rect 10672 4382 10678 4399
rect 10695 4382 10701 4399
rect 10672 4365 10701 4382
rect 10672 4348 10678 4365
rect 10695 4348 10701 4365
rect 10672 4340 10701 4348
rect 10716 4340 10737 4440
rect 10752 4433 10781 4440
rect 10752 4416 10758 4433
rect 10775 4416 10781 4433
rect 10752 4399 10781 4416
rect 10752 4382 10758 4399
rect 10775 4382 10781 4399
rect 10752 4365 10781 4382
rect 10752 4348 10758 4365
rect 10775 4348 10781 4365
rect 10752 4340 10781 4348
rect 10796 4433 10825 4440
rect 10796 4416 10802 4433
rect 10819 4416 10825 4433
rect 10796 4399 10825 4416
rect 10796 4382 10802 4399
rect 10819 4382 10825 4399
rect 10796 4365 10825 4382
rect 10796 4348 10802 4365
rect 10819 4348 10825 4365
rect 10796 4340 10825 4348
rect 10840 4433 10869 4440
rect 10840 4416 10846 4433
rect 10863 4416 10869 4433
rect 10840 4399 10869 4416
rect 10840 4382 10846 4399
rect 10863 4382 10869 4399
rect 10840 4365 10869 4382
rect 10840 4348 10846 4365
rect 10863 4348 10869 4365
rect 10840 4340 10869 4348
rect 10884 4340 10905 4440
rect 10920 4433 10949 4440
rect 10920 4416 10926 4433
rect 10943 4416 10949 4433
rect 10920 4399 10949 4416
rect 10920 4382 10926 4399
rect 10943 4382 10949 4399
rect 10920 4365 10949 4382
rect 10920 4348 10926 4365
rect 10943 4348 10949 4365
rect 10920 4340 10949 4348
rect 11250 4433 11279 4440
rect 11250 4416 11256 4433
rect 11273 4416 11279 4433
rect 11250 4399 11279 4416
rect 11250 4382 11256 4399
rect 11273 4382 11279 4399
rect 11250 4365 11279 4382
rect 11250 4348 11256 4365
rect 11273 4348 11279 4365
rect 11250 4340 11279 4348
rect 11294 4340 11315 4440
rect 11330 4433 11359 4440
rect 11330 4416 11336 4433
rect 11353 4416 11359 4433
rect 11330 4399 11359 4416
rect 11330 4382 11336 4399
rect 11353 4382 11359 4399
rect 11330 4365 11359 4382
rect 11330 4348 11336 4365
rect 11353 4348 11359 4365
rect 11330 4340 11359 4348
rect 11374 4433 11403 4440
rect 11374 4416 11380 4433
rect 11397 4416 11403 4433
rect 11374 4399 11403 4416
rect 11374 4382 11380 4399
rect 11397 4382 11403 4399
rect 11374 4365 11403 4382
rect 11374 4348 11380 4365
rect 11397 4348 11403 4365
rect 11374 4340 11403 4348
rect 11418 4433 11447 4440
rect 11418 4416 11424 4433
rect 11441 4416 11447 4433
rect 11418 4399 11447 4416
rect 11418 4382 11424 4399
rect 11441 4382 11447 4399
rect 11418 4365 11447 4382
rect 11418 4348 11424 4365
rect 11441 4348 11447 4365
rect 11418 4340 11447 4348
rect 11462 4340 11483 4440
rect 11498 4433 11527 4440
rect 11498 4416 11504 4433
rect 11521 4416 11527 4433
rect 11498 4399 11527 4416
rect 11498 4382 11504 4399
rect 11521 4382 11527 4399
rect 11498 4365 11527 4382
rect 11498 4348 11504 4365
rect 11521 4348 11527 4365
rect 11498 4340 11527 4348
rect 11861 4433 11890 4440
rect 11861 4416 11867 4433
rect 11884 4416 11890 4433
rect 11861 4399 11890 4416
rect 11861 4382 11867 4399
rect 11884 4382 11890 4399
rect 11861 4365 11890 4382
rect 11861 4348 11867 4365
rect 11884 4348 11890 4365
rect 11861 4340 11890 4348
rect 11905 4340 11926 4440
rect 11941 4433 11970 4440
rect 11941 4416 11947 4433
rect 11964 4416 11970 4433
rect 11941 4399 11970 4416
rect 11941 4382 11947 4399
rect 11964 4382 11970 4399
rect 11941 4365 11970 4382
rect 11941 4348 11947 4365
rect 11964 4348 11970 4365
rect 11941 4340 11970 4348
rect 11985 4433 12014 4440
rect 11985 4416 11991 4433
rect 12008 4416 12014 4433
rect 11985 4399 12014 4416
rect 11985 4382 11991 4399
rect 12008 4382 12014 4399
rect 11985 4365 12014 4382
rect 11985 4348 11991 4365
rect 12008 4348 12014 4365
rect 11985 4340 12014 4348
rect 12029 4433 12058 4440
rect 12029 4416 12035 4433
rect 12052 4416 12058 4433
rect 12029 4399 12058 4416
rect 12029 4382 12035 4399
rect 12052 4382 12058 4399
rect 12029 4365 12058 4382
rect 12029 4348 12035 4365
rect 12052 4348 12058 4365
rect 12029 4340 12058 4348
rect 12073 4340 12094 4440
rect 12109 4433 12138 4440
rect 12109 4416 12115 4433
rect 12132 4416 12138 4433
rect 12109 4399 12138 4416
rect 12109 4382 12115 4399
rect 12132 4382 12138 4399
rect 12109 4365 12138 4382
rect 12109 4348 12115 4365
rect 12132 4348 12138 4365
rect 12109 4340 12138 4348
rect 12472 4433 12501 4440
rect 12472 4416 12478 4433
rect 12495 4416 12501 4433
rect 12472 4399 12501 4416
rect 12472 4382 12478 4399
rect 12495 4382 12501 4399
rect 12472 4365 12501 4382
rect 12472 4348 12478 4365
rect 12495 4348 12501 4365
rect 12472 4340 12501 4348
rect 12516 4340 12537 4440
rect 12552 4433 12581 4440
rect 12552 4416 12558 4433
rect 12575 4416 12581 4433
rect 12552 4399 12581 4416
rect 12552 4382 12558 4399
rect 12575 4382 12581 4399
rect 12552 4365 12581 4382
rect 12552 4348 12558 4365
rect 12575 4348 12581 4365
rect 12552 4340 12581 4348
rect 12596 4433 12625 4440
rect 12596 4416 12602 4433
rect 12619 4416 12625 4433
rect 12596 4399 12625 4416
rect 12596 4382 12602 4399
rect 12619 4382 12625 4399
rect 12596 4365 12625 4382
rect 12596 4348 12602 4365
rect 12619 4348 12625 4365
rect 12596 4340 12625 4348
rect 12640 4433 12669 4440
rect 12640 4416 12646 4433
rect 12663 4416 12669 4433
rect 12640 4399 12669 4416
rect 12640 4382 12646 4399
rect 12663 4382 12669 4399
rect 12640 4365 12669 4382
rect 12640 4348 12646 4365
rect 12663 4348 12669 4365
rect 12640 4340 12669 4348
rect 12684 4340 12705 4440
rect 12720 4433 12749 4440
rect 12720 4416 12726 4433
rect 12743 4416 12749 4433
rect 12720 4399 12749 4416
rect 12720 4382 12726 4399
rect 12743 4382 12749 4399
rect 12720 4365 12749 4382
rect 12720 4348 12726 4365
rect 12743 4348 12749 4365
rect 12720 4340 12749 4348
<< pdiff >>
rect 10141 8039 10170 8044
rect 10141 8022 10147 8039
rect 10164 8022 10170 8039
rect 10141 8005 10170 8022
rect 10141 7988 10147 8005
rect 10164 7988 10170 8005
rect 10141 7971 10170 7988
rect 10141 7954 10147 7971
rect 10164 7954 10170 7971
rect 10141 7937 10170 7954
rect 10141 7920 10147 7937
rect 10164 7920 10170 7937
rect 10141 7903 10170 7920
rect 10141 7886 10147 7903
rect 10164 7886 10170 7903
rect 10141 7869 10170 7886
rect 10141 7852 10147 7869
rect 10164 7852 10170 7869
rect 10141 7844 10170 7852
rect 10185 8039 10214 8044
rect 10185 8022 10191 8039
rect 10208 8022 10214 8039
rect 10185 8005 10214 8022
rect 10185 7988 10191 8005
rect 10208 7988 10214 8005
rect 10185 7971 10214 7988
rect 10185 7954 10191 7971
rect 10208 7954 10214 7971
rect 10185 7937 10214 7954
rect 10185 7920 10191 7937
rect 10208 7920 10214 7937
rect 10185 7903 10214 7920
rect 10185 7886 10191 7903
rect 10208 7886 10214 7903
rect 10185 7869 10214 7886
rect 10185 7852 10191 7869
rect 10208 7852 10214 7869
rect 10185 7844 10214 7852
rect 10229 8039 10258 8044
rect 10229 8022 10235 8039
rect 10252 8022 10258 8039
rect 10229 8005 10258 8022
rect 10229 7988 10235 8005
rect 10252 7988 10258 8005
rect 10229 7971 10258 7988
rect 10229 7954 10235 7971
rect 10252 7954 10258 7971
rect 10229 7937 10258 7954
rect 10229 7920 10235 7937
rect 10252 7920 10258 7937
rect 10229 7903 10258 7920
rect 10229 7886 10235 7903
rect 10252 7886 10258 7903
rect 10229 7869 10258 7886
rect 10229 7852 10235 7869
rect 10252 7852 10258 7869
rect 10229 7844 10258 7852
rect 10752 8039 10781 8044
rect 10752 8022 10758 8039
rect 10775 8022 10781 8039
rect 10752 8005 10781 8022
rect 10752 7988 10758 8005
rect 10775 7988 10781 8005
rect 10752 7971 10781 7988
rect 10752 7954 10758 7971
rect 10775 7954 10781 7971
rect 10752 7937 10781 7954
rect 10752 7920 10758 7937
rect 10775 7920 10781 7937
rect 10752 7903 10781 7920
rect 10752 7886 10758 7903
rect 10775 7886 10781 7903
rect 10752 7869 10781 7886
rect 10752 7852 10758 7869
rect 10775 7852 10781 7869
rect 10752 7844 10781 7852
rect 10796 8039 10825 8044
rect 10796 8022 10802 8039
rect 10819 8022 10825 8039
rect 10796 8005 10825 8022
rect 10796 7988 10802 8005
rect 10819 7988 10825 8005
rect 10796 7971 10825 7988
rect 10796 7954 10802 7971
rect 10819 7954 10825 7971
rect 10796 7937 10825 7954
rect 10796 7920 10802 7937
rect 10819 7920 10825 7937
rect 10796 7903 10825 7920
rect 10796 7886 10802 7903
rect 10819 7886 10825 7903
rect 10796 7869 10825 7886
rect 10796 7852 10802 7869
rect 10819 7852 10825 7869
rect 10796 7844 10825 7852
rect 10840 8039 10869 8044
rect 10840 8022 10846 8039
rect 10863 8022 10869 8039
rect 10840 8005 10869 8022
rect 10840 7988 10846 8005
rect 10863 7988 10869 8005
rect 10840 7971 10869 7988
rect 10840 7954 10846 7971
rect 10863 7954 10869 7971
rect 10840 7937 10869 7954
rect 10840 7920 10846 7937
rect 10863 7920 10869 7937
rect 10840 7903 10869 7920
rect 10840 7886 10846 7903
rect 10863 7886 10869 7903
rect 10840 7869 10869 7886
rect 10840 7852 10846 7869
rect 10863 7852 10869 7869
rect 10840 7844 10869 7852
rect 11330 8039 11359 8044
rect 11330 8022 11336 8039
rect 11353 8022 11359 8039
rect 11330 8005 11359 8022
rect 11330 7988 11336 8005
rect 11353 7988 11359 8005
rect 11330 7971 11359 7988
rect 11330 7954 11336 7971
rect 11353 7954 11359 7971
rect 11330 7937 11359 7954
rect 11330 7920 11336 7937
rect 11353 7920 11359 7937
rect 11330 7903 11359 7920
rect 11330 7886 11336 7903
rect 11353 7886 11359 7903
rect 11330 7869 11359 7886
rect 11330 7852 11336 7869
rect 11353 7852 11359 7869
rect 11330 7844 11359 7852
rect 11374 8039 11403 8044
rect 11374 8022 11380 8039
rect 11397 8022 11403 8039
rect 11374 8005 11403 8022
rect 11374 7988 11380 8005
rect 11397 7988 11403 8005
rect 11374 7971 11403 7988
rect 11374 7954 11380 7971
rect 11397 7954 11403 7971
rect 11374 7937 11403 7954
rect 11374 7920 11380 7937
rect 11397 7920 11403 7937
rect 11374 7903 11403 7920
rect 11374 7886 11380 7903
rect 11397 7886 11403 7903
rect 11374 7869 11403 7886
rect 11374 7852 11380 7869
rect 11397 7852 11403 7869
rect 11374 7844 11403 7852
rect 11418 8039 11447 8044
rect 11418 8022 11424 8039
rect 11441 8022 11447 8039
rect 11418 8005 11447 8022
rect 11418 7988 11424 8005
rect 11441 7988 11447 8005
rect 11418 7971 11447 7988
rect 11418 7954 11424 7971
rect 11441 7954 11447 7971
rect 11418 7937 11447 7954
rect 11418 7920 11424 7937
rect 11441 7920 11447 7937
rect 11418 7903 11447 7920
rect 11418 7886 11424 7903
rect 11441 7886 11447 7903
rect 11418 7869 11447 7886
rect 11418 7852 11424 7869
rect 11441 7852 11447 7869
rect 11418 7844 11447 7852
rect 11941 8039 11970 8044
rect 11941 8022 11947 8039
rect 11964 8022 11970 8039
rect 11941 8005 11970 8022
rect 11941 7988 11947 8005
rect 11964 7988 11970 8005
rect 11941 7971 11970 7988
rect 11941 7954 11947 7971
rect 11964 7954 11970 7971
rect 11941 7937 11970 7954
rect 11941 7920 11947 7937
rect 11964 7920 11970 7937
rect 11941 7903 11970 7920
rect 11941 7886 11947 7903
rect 11964 7886 11970 7903
rect 11941 7869 11970 7886
rect 11941 7852 11947 7869
rect 11964 7852 11970 7869
rect 11941 7844 11970 7852
rect 11985 8039 12014 8044
rect 11985 8022 11991 8039
rect 12008 8022 12014 8039
rect 11985 8005 12014 8022
rect 11985 7988 11991 8005
rect 12008 7988 12014 8005
rect 11985 7971 12014 7988
rect 11985 7954 11991 7971
rect 12008 7954 12014 7971
rect 11985 7937 12014 7954
rect 11985 7920 11991 7937
rect 12008 7920 12014 7937
rect 11985 7903 12014 7920
rect 11985 7886 11991 7903
rect 12008 7886 12014 7903
rect 11985 7869 12014 7886
rect 11985 7852 11991 7869
rect 12008 7852 12014 7869
rect 11985 7844 12014 7852
rect 12029 8039 12058 8044
rect 12029 8022 12035 8039
rect 12052 8022 12058 8039
rect 12029 8005 12058 8022
rect 12029 7988 12035 8005
rect 12052 7988 12058 8005
rect 12029 7971 12058 7988
rect 12029 7954 12035 7971
rect 12052 7954 12058 7971
rect 12029 7937 12058 7954
rect 12029 7920 12035 7937
rect 12052 7920 12058 7937
rect 12029 7903 12058 7920
rect 12029 7886 12035 7903
rect 12052 7886 12058 7903
rect 12029 7869 12058 7886
rect 12029 7852 12035 7869
rect 12052 7852 12058 7869
rect 12029 7844 12058 7852
rect 12552 8039 12581 8044
rect 12552 8022 12558 8039
rect 12575 8022 12581 8039
rect 12552 8005 12581 8022
rect 12552 7988 12558 8005
rect 12575 7988 12581 8005
rect 12552 7971 12581 7988
rect 12552 7954 12558 7971
rect 12575 7954 12581 7971
rect 12552 7937 12581 7954
rect 12552 7920 12558 7937
rect 12575 7920 12581 7937
rect 12552 7903 12581 7920
rect 12552 7886 12558 7903
rect 12575 7886 12581 7903
rect 12552 7869 12581 7886
rect 12552 7852 12558 7869
rect 12575 7852 12581 7869
rect 12552 7844 12581 7852
rect 12596 8039 12625 8044
rect 12596 8022 12602 8039
rect 12619 8022 12625 8039
rect 12596 8005 12625 8022
rect 12596 7988 12602 8005
rect 12619 7988 12625 8005
rect 12596 7971 12625 7988
rect 12596 7954 12602 7971
rect 12619 7954 12625 7971
rect 12596 7937 12625 7954
rect 12596 7920 12602 7937
rect 12619 7920 12625 7937
rect 12596 7903 12625 7920
rect 12596 7886 12602 7903
rect 12619 7886 12625 7903
rect 12596 7869 12625 7886
rect 12596 7852 12602 7869
rect 12619 7852 12625 7869
rect 12596 7844 12625 7852
rect 12640 8039 12669 8044
rect 12640 8022 12646 8039
rect 12663 8022 12669 8039
rect 12640 8005 12669 8022
rect 12640 7988 12646 8005
rect 12663 7988 12669 8005
rect 12640 7971 12669 7988
rect 12640 7954 12646 7971
rect 12663 7954 12669 7971
rect 12640 7937 12669 7954
rect 12640 7920 12646 7937
rect 12663 7920 12669 7937
rect 12640 7903 12669 7920
rect 12640 7886 12646 7903
rect 12663 7886 12669 7903
rect 12640 7869 12669 7886
rect 12640 7852 12646 7869
rect 12663 7852 12669 7869
rect 12640 7844 12669 7852
rect 9530 7389 9559 7394
rect 9530 7372 9536 7389
rect 9553 7372 9559 7389
rect 9530 7355 9559 7372
rect 9530 7338 9536 7355
rect 9553 7338 9559 7355
rect 9530 7321 9559 7338
rect 9530 7304 9536 7321
rect 9553 7304 9559 7321
rect 9530 7287 9559 7304
rect 9530 7270 9536 7287
rect 9553 7270 9559 7287
rect 9530 7253 9559 7270
rect 9530 7236 9536 7253
rect 9553 7236 9559 7253
rect 9530 7219 9559 7236
rect 9530 7202 9536 7219
rect 9553 7202 9559 7219
rect 9530 7194 9559 7202
rect 9574 7389 9603 7394
rect 9574 7372 9580 7389
rect 9597 7372 9603 7389
rect 9574 7355 9603 7372
rect 9574 7338 9580 7355
rect 9597 7338 9603 7355
rect 9574 7321 9603 7338
rect 9574 7304 9580 7321
rect 9597 7304 9603 7321
rect 9574 7287 9603 7304
rect 9574 7270 9580 7287
rect 9597 7270 9603 7287
rect 9574 7253 9603 7270
rect 9574 7236 9580 7253
rect 9597 7236 9603 7253
rect 9574 7219 9603 7236
rect 9574 7202 9580 7219
rect 9597 7202 9603 7219
rect 9574 7194 9603 7202
rect 9618 7389 9647 7394
rect 9618 7372 9624 7389
rect 9641 7372 9647 7389
rect 9618 7355 9647 7372
rect 9618 7338 9624 7355
rect 9641 7338 9647 7355
rect 9618 7321 9647 7338
rect 9618 7304 9624 7321
rect 9641 7304 9647 7321
rect 9618 7287 9647 7304
rect 9618 7270 9624 7287
rect 9641 7270 9647 7287
rect 9618 7253 9647 7270
rect 9618 7236 9624 7253
rect 9641 7236 9647 7253
rect 9618 7219 9647 7236
rect 9618 7202 9624 7219
rect 9641 7202 9647 7219
rect 9618 7194 9647 7202
rect 10141 7389 10170 7394
rect 10141 7372 10147 7389
rect 10164 7372 10170 7389
rect 10141 7355 10170 7372
rect 10141 7338 10147 7355
rect 10164 7338 10170 7355
rect 10141 7321 10170 7338
rect 10141 7304 10147 7321
rect 10164 7304 10170 7321
rect 10141 7287 10170 7304
rect 10141 7270 10147 7287
rect 10164 7270 10170 7287
rect 10141 7253 10170 7270
rect 10141 7236 10147 7253
rect 10164 7236 10170 7253
rect 10141 7219 10170 7236
rect 10141 7202 10147 7219
rect 10164 7202 10170 7219
rect 10141 7194 10170 7202
rect 10185 7389 10214 7394
rect 10185 7372 10191 7389
rect 10208 7372 10214 7389
rect 10185 7355 10214 7372
rect 10185 7338 10191 7355
rect 10208 7338 10214 7355
rect 10185 7321 10214 7338
rect 10185 7304 10191 7321
rect 10208 7304 10214 7321
rect 10185 7287 10214 7304
rect 10185 7270 10191 7287
rect 10208 7270 10214 7287
rect 10185 7253 10214 7270
rect 10185 7236 10191 7253
rect 10208 7236 10214 7253
rect 10185 7219 10214 7236
rect 10185 7202 10191 7219
rect 10208 7202 10214 7219
rect 10185 7194 10214 7202
rect 10229 7389 10258 7394
rect 10229 7372 10235 7389
rect 10252 7372 10258 7389
rect 10229 7355 10258 7372
rect 10229 7338 10235 7355
rect 10252 7338 10258 7355
rect 10229 7321 10258 7338
rect 10229 7304 10235 7321
rect 10252 7304 10258 7321
rect 10229 7287 10258 7304
rect 10229 7270 10235 7287
rect 10252 7270 10258 7287
rect 10229 7253 10258 7270
rect 10229 7236 10235 7253
rect 10252 7236 10258 7253
rect 10229 7219 10258 7236
rect 10229 7202 10235 7219
rect 10252 7202 10258 7219
rect 10229 7194 10258 7202
rect 10752 7389 10781 7394
rect 10752 7372 10758 7389
rect 10775 7372 10781 7389
rect 10752 7355 10781 7372
rect 10752 7338 10758 7355
rect 10775 7338 10781 7355
rect 10752 7321 10781 7338
rect 10752 7304 10758 7321
rect 10775 7304 10781 7321
rect 10752 7287 10781 7304
rect 10752 7270 10758 7287
rect 10775 7270 10781 7287
rect 10752 7253 10781 7270
rect 10752 7236 10758 7253
rect 10775 7236 10781 7253
rect 10752 7219 10781 7236
rect 10752 7202 10758 7219
rect 10775 7202 10781 7219
rect 10752 7194 10781 7202
rect 10796 7389 10825 7394
rect 10796 7372 10802 7389
rect 10819 7372 10825 7389
rect 10796 7355 10825 7372
rect 10796 7338 10802 7355
rect 10819 7338 10825 7355
rect 10796 7321 10825 7338
rect 10796 7304 10802 7321
rect 10819 7304 10825 7321
rect 10796 7287 10825 7304
rect 10796 7270 10802 7287
rect 10819 7270 10825 7287
rect 10796 7253 10825 7270
rect 10796 7236 10802 7253
rect 10819 7236 10825 7253
rect 10796 7219 10825 7236
rect 10796 7202 10802 7219
rect 10819 7202 10825 7219
rect 10796 7194 10825 7202
rect 10840 7389 10869 7394
rect 10840 7372 10846 7389
rect 10863 7372 10869 7389
rect 10840 7355 10869 7372
rect 10840 7338 10846 7355
rect 10863 7338 10869 7355
rect 10840 7321 10869 7338
rect 10840 7304 10846 7321
rect 10863 7304 10869 7321
rect 10840 7287 10869 7304
rect 10840 7270 10846 7287
rect 10863 7270 10869 7287
rect 10840 7253 10869 7270
rect 10840 7236 10846 7253
rect 10863 7236 10869 7253
rect 10840 7219 10869 7236
rect 10840 7202 10846 7219
rect 10863 7202 10869 7219
rect 10840 7194 10869 7202
rect 11330 7389 11359 7394
rect 11330 7372 11336 7389
rect 11353 7372 11359 7389
rect 11330 7355 11359 7372
rect 11330 7338 11336 7355
rect 11353 7338 11359 7355
rect 11330 7321 11359 7338
rect 11330 7304 11336 7321
rect 11353 7304 11359 7321
rect 11330 7287 11359 7304
rect 11330 7270 11336 7287
rect 11353 7270 11359 7287
rect 11330 7253 11359 7270
rect 11330 7236 11336 7253
rect 11353 7236 11359 7253
rect 11330 7219 11359 7236
rect 11330 7202 11336 7219
rect 11353 7202 11359 7219
rect 11330 7194 11359 7202
rect 11374 7389 11403 7394
rect 11374 7372 11380 7389
rect 11397 7372 11403 7389
rect 11374 7355 11403 7372
rect 11374 7338 11380 7355
rect 11397 7338 11403 7355
rect 11374 7321 11403 7338
rect 11374 7304 11380 7321
rect 11397 7304 11403 7321
rect 11374 7287 11403 7304
rect 11374 7270 11380 7287
rect 11397 7270 11403 7287
rect 11374 7253 11403 7270
rect 11374 7236 11380 7253
rect 11397 7236 11403 7253
rect 11374 7219 11403 7236
rect 11374 7202 11380 7219
rect 11397 7202 11403 7219
rect 11374 7194 11403 7202
rect 11418 7389 11447 7394
rect 11418 7372 11424 7389
rect 11441 7372 11447 7389
rect 11418 7355 11447 7372
rect 11418 7338 11424 7355
rect 11441 7338 11447 7355
rect 11418 7321 11447 7338
rect 11418 7304 11424 7321
rect 11441 7304 11447 7321
rect 11418 7287 11447 7304
rect 11418 7270 11424 7287
rect 11441 7270 11447 7287
rect 11418 7253 11447 7270
rect 11418 7236 11424 7253
rect 11441 7236 11447 7253
rect 11418 7219 11447 7236
rect 11418 7202 11424 7219
rect 11441 7202 11447 7219
rect 11418 7194 11447 7202
rect 11941 7389 11970 7394
rect 11941 7372 11947 7389
rect 11964 7372 11970 7389
rect 11941 7355 11970 7372
rect 11941 7338 11947 7355
rect 11964 7338 11970 7355
rect 11941 7321 11970 7338
rect 11941 7304 11947 7321
rect 11964 7304 11970 7321
rect 11941 7287 11970 7304
rect 11941 7270 11947 7287
rect 11964 7270 11970 7287
rect 11941 7253 11970 7270
rect 11941 7236 11947 7253
rect 11964 7236 11970 7253
rect 11941 7219 11970 7236
rect 11941 7202 11947 7219
rect 11964 7202 11970 7219
rect 11941 7194 11970 7202
rect 11985 7389 12014 7394
rect 11985 7372 11991 7389
rect 12008 7372 12014 7389
rect 11985 7355 12014 7372
rect 11985 7338 11991 7355
rect 12008 7338 12014 7355
rect 11985 7321 12014 7338
rect 11985 7304 11991 7321
rect 12008 7304 12014 7321
rect 11985 7287 12014 7304
rect 11985 7270 11991 7287
rect 12008 7270 12014 7287
rect 11985 7253 12014 7270
rect 11985 7236 11991 7253
rect 12008 7236 12014 7253
rect 11985 7219 12014 7236
rect 11985 7202 11991 7219
rect 12008 7202 12014 7219
rect 11985 7194 12014 7202
rect 12029 7389 12058 7394
rect 12029 7372 12035 7389
rect 12052 7372 12058 7389
rect 12029 7355 12058 7372
rect 12029 7338 12035 7355
rect 12052 7338 12058 7355
rect 12029 7321 12058 7338
rect 12029 7304 12035 7321
rect 12052 7304 12058 7321
rect 12029 7287 12058 7304
rect 12029 7270 12035 7287
rect 12052 7270 12058 7287
rect 12029 7253 12058 7270
rect 12029 7236 12035 7253
rect 12052 7236 12058 7253
rect 12029 7219 12058 7236
rect 12029 7202 12035 7219
rect 12052 7202 12058 7219
rect 12029 7194 12058 7202
rect 12552 7389 12581 7394
rect 12552 7372 12558 7389
rect 12575 7372 12581 7389
rect 12552 7355 12581 7372
rect 12552 7338 12558 7355
rect 12575 7338 12581 7355
rect 12552 7321 12581 7338
rect 12552 7304 12558 7321
rect 12575 7304 12581 7321
rect 12552 7287 12581 7304
rect 12552 7270 12558 7287
rect 12575 7270 12581 7287
rect 12552 7253 12581 7270
rect 12552 7236 12558 7253
rect 12575 7236 12581 7253
rect 12552 7219 12581 7236
rect 12552 7202 12558 7219
rect 12575 7202 12581 7219
rect 12552 7194 12581 7202
rect 12596 7389 12625 7394
rect 12596 7372 12602 7389
rect 12619 7372 12625 7389
rect 12596 7355 12625 7372
rect 12596 7338 12602 7355
rect 12619 7338 12625 7355
rect 12596 7321 12625 7338
rect 12596 7304 12602 7321
rect 12619 7304 12625 7321
rect 12596 7287 12625 7304
rect 12596 7270 12602 7287
rect 12619 7270 12625 7287
rect 12596 7253 12625 7270
rect 12596 7236 12602 7253
rect 12619 7236 12625 7253
rect 12596 7219 12625 7236
rect 12596 7202 12602 7219
rect 12619 7202 12625 7219
rect 12596 7194 12625 7202
rect 12640 7389 12669 7394
rect 12640 7372 12646 7389
rect 12663 7372 12669 7389
rect 12640 7355 12669 7372
rect 12640 7338 12646 7355
rect 12663 7338 12669 7355
rect 12640 7321 12669 7338
rect 12640 7304 12646 7321
rect 12663 7304 12669 7321
rect 12640 7287 12669 7304
rect 12640 7270 12646 7287
rect 12663 7270 12669 7287
rect 12640 7253 12669 7270
rect 12640 7236 12646 7253
rect 12663 7236 12669 7253
rect 12640 7219 12669 7236
rect 12640 7202 12646 7219
rect 12663 7202 12669 7219
rect 12640 7194 12669 7202
rect 9530 6749 9559 6754
rect 9530 6732 9536 6749
rect 9553 6732 9559 6749
rect 9530 6715 9559 6732
rect 9530 6698 9536 6715
rect 9553 6698 9559 6715
rect 9530 6681 9559 6698
rect 9530 6664 9536 6681
rect 9553 6664 9559 6681
rect 9530 6647 9559 6664
rect 9530 6630 9536 6647
rect 9553 6630 9559 6647
rect 9530 6613 9559 6630
rect 9530 6596 9536 6613
rect 9553 6596 9559 6613
rect 9530 6579 9559 6596
rect 9530 6562 9536 6579
rect 9553 6562 9559 6579
rect 9530 6554 9559 6562
rect 9574 6749 9603 6754
rect 9574 6732 9580 6749
rect 9597 6732 9603 6749
rect 9574 6715 9603 6732
rect 9574 6698 9580 6715
rect 9597 6698 9603 6715
rect 9574 6681 9603 6698
rect 9574 6664 9580 6681
rect 9597 6664 9603 6681
rect 9574 6647 9603 6664
rect 9574 6630 9580 6647
rect 9597 6630 9603 6647
rect 9574 6613 9603 6630
rect 9574 6596 9580 6613
rect 9597 6596 9603 6613
rect 9574 6579 9603 6596
rect 9574 6562 9580 6579
rect 9597 6562 9603 6579
rect 9574 6554 9603 6562
rect 9618 6749 9647 6754
rect 9618 6732 9624 6749
rect 9641 6732 9647 6749
rect 9618 6715 9647 6732
rect 9618 6698 9624 6715
rect 9641 6698 9647 6715
rect 9618 6681 9647 6698
rect 9618 6664 9624 6681
rect 9641 6664 9647 6681
rect 9618 6647 9647 6664
rect 9618 6630 9624 6647
rect 9641 6630 9647 6647
rect 9618 6613 9647 6630
rect 9618 6596 9624 6613
rect 9641 6596 9647 6613
rect 9618 6579 9647 6596
rect 9618 6562 9624 6579
rect 9641 6562 9647 6579
rect 9618 6554 9647 6562
rect 10141 6749 10170 6754
rect 10141 6732 10147 6749
rect 10164 6732 10170 6749
rect 10141 6715 10170 6732
rect 10141 6698 10147 6715
rect 10164 6698 10170 6715
rect 10141 6681 10170 6698
rect 10141 6664 10147 6681
rect 10164 6664 10170 6681
rect 10141 6647 10170 6664
rect 10141 6630 10147 6647
rect 10164 6630 10170 6647
rect 10141 6613 10170 6630
rect 10141 6596 10147 6613
rect 10164 6596 10170 6613
rect 10141 6579 10170 6596
rect 10141 6562 10147 6579
rect 10164 6562 10170 6579
rect 10141 6554 10170 6562
rect 10185 6749 10214 6754
rect 10185 6732 10191 6749
rect 10208 6732 10214 6749
rect 10185 6715 10214 6732
rect 10185 6698 10191 6715
rect 10208 6698 10214 6715
rect 10185 6681 10214 6698
rect 10185 6664 10191 6681
rect 10208 6664 10214 6681
rect 10185 6647 10214 6664
rect 10185 6630 10191 6647
rect 10208 6630 10214 6647
rect 10185 6613 10214 6630
rect 10185 6596 10191 6613
rect 10208 6596 10214 6613
rect 10185 6579 10214 6596
rect 10185 6562 10191 6579
rect 10208 6562 10214 6579
rect 10185 6554 10214 6562
rect 10229 6749 10258 6754
rect 10229 6732 10235 6749
rect 10252 6732 10258 6749
rect 10229 6715 10258 6732
rect 10229 6698 10235 6715
rect 10252 6698 10258 6715
rect 10229 6681 10258 6698
rect 10229 6664 10235 6681
rect 10252 6664 10258 6681
rect 10229 6647 10258 6664
rect 10229 6630 10235 6647
rect 10252 6630 10258 6647
rect 10229 6613 10258 6630
rect 10229 6596 10235 6613
rect 10252 6596 10258 6613
rect 10229 6579 10258 6596
rect 10229 6562 10235 6579
rect 10252 6562 10258 6579
rect 10229 6554 10258 6562
rect 10752 6749 10781 6754
rect 10752 6732 10758 6749
rect 10775 6732 10781 6749
rect 10752 6715 10781 6732
rect 10752 6698 10758 6715
rect 10775 6698 10781 6715
rect 10752 6681 10781 6698
rect 10752 6664 10758 6681
rect 10775 6664 10781 6681
rect 10752 6647 10781 6664
rect 10752 6630 10758 6647
rect 10775 6630 10781 6647
rect 10752 6613 10781 6630
rect 10752 6596 10758 6613
rect 10775 6596 10781 6613
rect 10752 6579 10781 6596
rect 10752 6562 10758 6579
rect 10775 6562 10781 6579
rect 10752 6554 10781 6562
rect 10796 6749 10825 6754
rect 10796 6732 10802 6749
rect 10819 6732 10825 6749
rect 10796 6715 10825 6732
rect 10796 6698 10802 6715
rect 10819 6698 10825 6715
rect 10796 6681 10825 6698
rect 10796 6664 10802 6681
rect 10819 6664 10825 6681
rect 10796 6647 10825 6664
rect 10796 6630 10802 6647
rect 10819 6630 10825 6647
rect 10796 6613 10825 6630
rect 10796 6596 10802 6613
rect 10819 6596 10825 6613
rect 10796 6579 10825 6596
rect 10796 6562 10802 6579
rect 10819 6562 10825 6579
rect 10796 6554 10825 6562
rect 10840 6749 10869 6754
rect 10840 6732 10846 6749
rect 10863 6732 10869 6749
rect 10840 6715 10869 6732
rect 10840 6698 10846 6715
rect 10863 6698 10869 6715
rect 10840 6681 10869 6698
rect 10840 6664 10846 6681
rect 10863 6664 10869 6681
rect 10840 6647 10869 6664
rect 10840 6630 10846 6647
rect 10863 6630 10869 6647
rect 10840 6613 10869 6630
rect 10840 6596 10846 6613
rect 10863 6596 10869 6613
rect 10840 6579 10869 6596
rect 10840 6562 10846 6579
rect 10863 6562 10869 6579
rect 10840 6554 10869 6562
rect 11330 6749 11359 6754
rect 11330 6732 11336 6749
rect 11353 6732 11359 6749
rect 11330 6715 11359 6732
rect 11330 6698 11336 6715
rect 11353 6698 11359 6715
rect 11330 6681 11359 6698
rect 11330 6664 11336 6681
rect 11353 6664 11359 6681
rect 11330 6647 11359 6664
rect 11330 6630 11336 6647
rect 11353 6630 11359 6647
rect 11330 6613 11359 6630
rect 11330 6596 11336 6613
rect 11353 6596 11359 6613
rect 11330 6579 11359 6596
rect 11330 6562 11336 6579
rect 11353 6562 11359 6579
rect 11330 6554 11359 6562
rect 11374 6749 11403 6754
rect 11374 6732 11380 6749
rect 11397 6732 11403 6749
rect 11374 6715 11403 6732
rect 11374 6698 11380 6715
rect 11397 6698 11403 6715
rect 11374 6681 11403 6698
rect 11374 6664 11380 6681
rect 11397 6664 11403 6681
rect 11374 6647 11403 6664
rect 11374 6630 11380 6647
rect 11397 6630 11403 6647
rect 11374 6613 11403 6630
rect 11374 6596 11380 6613
rect 11397 6596 11403 6613
rect 11374 6579 11403 6596
rect 11374 6562 11380 6579
rect 11397 6562 11403 6579
rect 11374 6554 11403 6562
rect 11418 6749 11447 6754
rect 11418 6732 11424 6749
rect 11441 6732 11447 6749
rect 11418 6715 11447 6732
rect 11418 6698 11424 6715
rect 11441 6698 11447 6715
rect 11418 6681 11447 6698
rect 11418 6664 11424 6681
rect 11441 6664 11447 6681
rect 11418 6647 11447 6664
rect 11418 6630 11424 6647
rect 11441 6630 11447 6647
rect 11418 6613 11447 6630
rect 11418 6596 11424 6613
rect 11441 6596 11447 6613
rect 11418 6579 11447 6596
rect 11418 6562 11424 6579
rect 11441 6562 11447 6579
rect 11418 6554 11447 6562
rect 11941 6749 11970 6754
rect 11941 6732 11947 6749
rect 11964 6732 11970 6749
rect 11941 6715 11970 6732
rect 11941 6698 11947 6715
rect 11964 6698 11970 6715
rect 11941 6681 11970 6698
rect 11941 6664 11947 6681
rect 11964 6664 11970 6681
rect 11941 6647 11970 6664
rect 11941 6630 11947 6647
rect 11964 6630 11970 6647
rect 11941 6613 11970 6630
rect 11941 6596 11947 6613
rect 11964 6596 11970 6613
rect 11941 6579 11970 6596
rect 11941 6562 11947 6579
rect 11964 6562 11970 6579
rect 11941 6554 11970 6562
rect 11985 6749 12014 6754
rect 11985 6732 11991 6749
rect 12008 6732 12014 6749
rect 11985 6715 12014 6732
rect 11985 6698 11991 6715
rect 12008 6698 12014 6715
rect 11985 6681 12014 6698
rect 11985 6664 11991 6681
rect 12008 6664 12014 6681
rect 11985 6647 12014 6664
rect 11985 6630 11991 6647
rect 12008 6630 12014 6647
rect 11985 6613 12014 6630
rect 11985 6596 11991 6613
rect 12008 6596 12014 6613
rect 11985 6579 12014 6596
rect 11985 6562 11991 6579
rect 12008 6562 12014 6579
rect 11985 6554 12014 6562
rect 12029 6749 12058 6754
rect 12029 6732 12035 6749
rect 12052 6732 12058 6749
rect 12029 6715 12058 6732
rect 12029 6698 12035 6715
rect 12052 6698 12058 6715
rect 12029 6681 12058 6698
rect 12029 6664 12035 6681
rect 12052 6664 12058 6681
rect 12029 6647 12058 6664
rect 12029 6630 12035 6647
rect 12052 6630 12058 6647
rect 12029 6613 12058 6630
rect 12029 6596 12035 6613
rect 12052 6596 12058 6613
rect 12029 6579 12058 6596
rect 12029 6562 12035 6579
rect 12052 6562 12058 6579
rect 12029 6554 12058 6562
rect 12552 6749 12581 6754
rect 12552 6732 12558 6749
rect 12575 6732 12581 6749
rect 12552 6715 12581 6732
rect 12552 6698 12558 6715
rect 12575 6698 12581 6715
rect 12552 6681 12581 6698
rect 12552 6664 12558 6681
rect 12575 6664 12581 6681
rect 12552 6647 12581 6664
rect 12552 6630 12558 6647
rect 12575 6630 12581 6647
rect 12552 6613 12581 6630
rect 12552 6596 12558 6613
rect 12575 6596 12581 6613
rect 12552 6579 12581 6596
rect 12552 6562 12558 6579
rect 12575 6562 12581 6579
rect 12552 6554 12581 6562
rect 12596 6749 12625 6754
rect 12596 6732 12602 6749
rect 12619 6732 12625 6749
rect 12596 6715 12625 6732
rect 12596 6698 12602 6715
rect 12619 6698 12625 6715
rect 12596 6681 12625 6698
rect 12596 6664 12602 6681
rect 12619 6664 12625 6681
rect 12596 6647 12625 6664
rect 12596 6630 12602 6647
rect 12619 6630 12625 6647
rect 12596 6613 12625 6630
rect 12596 6596 12602 6613
rect 12619 6596 12625 6613
rect 12596 6579 12625 6596
rect 12596 6562 12602 6579
rect 12619 6562 12625 6579
rect 12596 6554 12625 6562
rect 12640 6749 12669 6754
rect 12640 6732 12646 6749
rect 12663 6732 12669 6749
rect 12640 6715 12669 6732
rect 12640 6698 12646 6715
rect 12663 6698 12669 6715
rect 12640 6681 12669 6698
rect 12640 6664 12646 6681
rect 12663 6664 12669 6681
rect 12640 6647 12669 6664
rect 12640 6630 12646 6647
rect 12663 6630 12669 6647
rect 12640 6613 12669 6630
rect 12640 6596 12646 6613
rect 12663 6596 12669 6613
rect 12640 6579 12669 6596
rect 12640 6562 12646 6579
rect 12663 6562 12669 6579
rect 12640 6554 12669 6562
rect 9530 6099 9559 6104
rect 9530 6082 9536 6099
rect 9553 6082 9559 6099
rect 9530 6065 9559 6082
rect 9530 6048 9536 6065
rect 9553 6048 9559 6065
rect 9530 6031 9559 6048
rect 9530 6014 9536 6031
rect 9553 6014 9559 6031
rect 9530 5997 9559 6014
rect 9530 5980 9536 5997
rect 9553 5980 9559 5997
rect 9530 5963 9559 5980
rect 9530 5946 9536 5963
rect 9553 5946 9559 5963
rect 9530 5929 9559 5946
rect 9530 5912 9536 5929
rect 9553 5912 9559 5929
rect 9530 5904 9559 5912
rect 9574 6099 9603 6104
rect 9574 6082 9580 6099
rect 9597 6082 9603 6099
rect 9574 6065 9603 6082
rect 9574 6048 9580 6065
rect 9597 6048 9603 6065
rect 9574 6031 9603 6048
rect 9574 6014 9580 6031
rect 9597 6014 9603 6031
rect 9574 5997 9603 6014
rect 9574 5980 9580 5997
rect 9597 5980 9603 5997
rect 9574 5963 9603 5980
rect 9574 5946 9580 5963
rect 9597 5946 9603 5963
rect 9574 5929 9603 5946
rect 9574 5912 9580 5929
rect 9597 5912 9603 5929
rect 9574 5904 9603 5912
rect 9618 6099 9647 6104
rect 9618 6082 9624 6099
rect 9641 6082 9647 6099
rect 9618 6065 9647 6082
rect 9618 6048 9624 6065
rect 9641 6048 9647 6065
rect 9618 6031 9647 6048
rect 9618 6014 9624 6031
rect 9641 6014 9647 6031
rect 9618 5997 9647 6014
rect 9618 5980 9624 5997
rect 9641 5980 9647 5997
rect 9618 5963 9647 5980
rect 9618 5946 9624 5963
rect 9641 5946 9647 5963
rect 9618 5929 9647 5946
rect 9618 5912 9624 5929
rect 9641 5912 9647 5929
rect 9618 5904 9647 5912
rect 10141 6099 10170 6104
rect 10141 6082 10147 6099
rect 10164 6082 10170 6099
rect 10141 6065 10170 6082
rect 10141 6048 10147 6065
rect 10164 6048 10170 6065
rect 10141 6031 10170 6048
rect 10141 6014 10147 6031
rect 10164 6014 10170 6031
rect 10141 5997 10170 6014
rect 10141 5980 10147 5997
rect 10164 5980 10170 5997
rect 10141 5963 10170 5980
rect 10141 5946 10147 5963
rect 10164 5946 10170 5963
rect 10141 5929 10170 5946
rect 10141 5912 10147 5929
rect 10164 5912 10170 5929
rect 10141 5904 10170 5912
rect 10185 6099 10214 6104
rect 10185 6082 10191 6099
rect 10208 6082 10214 6099
rect 10185 6065 10214 6082
rect 10185 6048 10191 6065
rect 10208 6048 10214 6065
rect 10185 6031 10214 6048
rect 10185 6014 10191 6031
rect 10208 6014 10214 6031
rect 10185 5997 10214 6014
rect 10185 5980 10191 5997
rect 10208 5980 10214 5997
rect 10185 5963 10214 5980
rect 10185 5946 10191 5963
rect 10208 5946 10214 5963
rect 10185 5929 10214 5946
rect 10185 5912 10191 5929
rect 10208 5912 10214 5929
rect 10185 5904 10214 5912
rect 10229 6099 10258 6104
rect 10229 6082 10235 6099
rect 10252 6082 10258 6099
rect 10229 6065 10258 6082
rect 10229 6048 10235 6065
rect 10252 6048 10258 6065
rect 10229 6031 10258 6048
rect 10229 6014 10235 6031
rect 10252 6014 10258 6031
rect 10229 5997 10258 6014
rect 10229 5980 10235 5997
rect 10252 5980 10258 5997
rect 10229 5963 10258 5980
rect 10229 5946 10235 5963
rect 10252 5946 10258 5963
rect 10229 5929 10258 5946
rect 10229 5912 10235 5929
rect 10252 5912 10258 5929
rect 10229 5904 10258 5912
rect 10752 6099 10781 6104
rect 10752 6082 10758 6099
rect 10775 6082 10781 6099
rect 10752 6065 10781 6082
rect 10752 6048 10758 6065
rect 10775 6048 10781 6065
rect 10752 6031 10781 6048
rect 10752 6014 10758 6031
rect 10775 6014 10781 6031
rect 10752 5997 10781 6014
rect 10752 5980 10758 5997
rect 10775 5980 10781 5997
rect 10752 5963 10781 5980
rect 10752 5946 10758 5963
rect 10775 5946 10781 5963
rect 10752 5929 10781 5946
rect 10752 5912 10758 5929
rect 10775 5912 10781 5929
rect 10752 5904 10781 5912
rect 10796 6099 10825 6104
rect 10796 6082 10802 6099
rect 10819 6082 10825 6099
rect 10796 6065 10825 6082
rect 10796 6048 10802 6065
rect 10819 6048 10825 6065
rect 10796 6031 10825 6048
rect 10796 6014 10802 6031
rect 10819 6014 10825 6031
rect 10796 5997 10825 6014
rect 10796 5980 10802 5997
rect 10819 5980 10825 5997
rect 10796 5963 10825 5980
rect 10796 5946 10802 5963
rect 10819 5946 10825 5963
rect 10796 5929 10825 5946
rect 10796 5912 10802 5929
rect 10819 5912 10825 5929
rect 10796 5904 10825 5912
rect 10840 6099 10869 6104
rect 10840 6082 10846 6099
rect 10863 6082 10869 6099
rect 10840 6065 10869 6082
rect 10840 6048 10846 6065
rect 10863 6048 10869 6065
rect 10840 6031 10869 6048
rect 10840 6014 10846 6031
rect 10863 6014 10869 6031
rect 10840 5997 10869 6014
rect 10840 5980 10846 5997
rect 10863 5980 10869 5997
rect 10840 5963 10869 5980
rect 10840 5946 10846 5963
rect 10863 5946 10869 5963
rect 10840 5929 10869 5946
rect 10840 5912 10846 5929
rect 10863 5912 10869 5929
rect 10840 5904 10869 5912
rect 11330 6099 11359 6104
rect 11330 6082 11336 6099
rect 11353 6082 11359 6099
rect 11330 6065 11359 6082
rect 11330 6048 11336 6065
rect 11353 6048 11359 6065
rect 11330 6031 11359 6048
rect 11330 6014 11336 6031
rect 11353 6014 11359 6031
rect 11330 5997 11359 6014
rect 11330 5980 11336 5997
rect 11353 5980 11359 5997
rect 11330 5963 11359 5980
rect 11330 5946 11336 5963
rect 11353 5946 11359 5963
rect 11330 5929 11359 5946
rect 11330 5912 11336 5929
rect 11353 5912 11359 5929
rect 11330 5904 11359 5912
rect 11374 6099 11403 6104
rect 11374 6082 11380 6099
rect 11397 6082 11403 6099
rect 11374 6065 11403 6082
rect 11374 6048 11380 6065
rect 11397 6048 11403 6065
rect 11374 6031 11403 6048
rect 11374 6014 11380 6031
rect 11397 6014 11403 6031
rect 11374 5997 11403 6014
rect 11374 5980 11380 5997
rect 11397 5980 11403 5997
rect 11374 5963 11403 5980
rect 11374 5946 11380 5963
rect 11397 5946 11403 5963
rect 11374 5929 11403 5946
rect 11374 5912 11380 5929
rect 11397 5912 11403 5929
rect 11374 5904 11403 5912
rect 11418 6099 11447 6104
rect 11418 6082 11424 6099
rect 11441 6082 11447 6099
rect 11418 6065 11447 6082
rect 11418 6048 11424 6065
rect 11441 6048 11447 6065
rect 11418 6031 11447 6048
rect 11418 6014 11424 6031
rect 11441 6014 11447 6031
rect 11418 5997 11447 6014
rect 11418 5980 11424 5997
rect 11441 5980 11447 5997
rect 11418 5963 11447 5980
rect 11418 5946 11424 5963
rect 11441 5946 11447 5963
rect 11418 5929 11447 5946
rect 11418 5912 11424 5929
rect 11441 5912 11447 5929
rect 11418 5904 11447 5912
rect 11941 6099 11970 6104
rect 11941 6082 11947 6099
rect 11964 6082 11970 6099
rect 11941 6065 11970 6082
rect 11941 6048 11947 6065
rect 11964 6048 11970 6065
rect 11941 6031 11970 6048
rect 11941 6014 11947 6031
rect 11964 6014 11970 6031
rect 11941 5997 11970 6014
rect 11941 5980 11947 5997
rect 11964 5980 11970 5997
rect 11941 5963 11970 5980
rect 11941 5946 11947 5963
rect 11964 5946 11970 5963
rect 11941 5929 11970 5946
rect 11941 5912 11947 5929
rect 11964 5912 11970 5929
rect 11941 5904 11970 5912
rect 11985 6099 12014 6104
rect 11985 6082 11991 6099
rect 12008 6082 12014 6099
rect 11985 6065 12014 6082
rect 11985 6048 11991 6065
rect 12008 6048 12014 6065
rect 11985 6031 12014 6048
rect 11985 6014 11991 6031
rect 12008 6014 12014 6031
rect 11985 5997 12014 6014
rect 11985 5980 11991 5997
rect 12008 5980 12014 5997
rect 11985 5963 12014 5980
rect 11985 5946 11991 5963
rect 12008 5946 12014 5963
rect 11985 5929 12014 5946
rect 11985 5912 11991 5929
rect 12008 5912 12014 5929
rect 11985 5904 12014 5912
rect 12029 6099 12058 6104
rect 12029 6082 12035 6099
rect 12052 6082 12058 6099
rect 12029 6065 12058 6082
rect 12029 6048 12035 6065
rect 12052 6048 12058 6065
rect 12029 6031 12058 6048
rect 12029 6014 12035 6031
rect 12052 6014 12058 6031
rect 12029 5997 12058 6014
rect 12029 5980 12035 5997
rect 12052 5980 12058 5997
rect 12029 5963 12058 5980
rect 12029 5946 12035 5963
rect 12052 5946 12058 5963
rect 12029 5929 12058 5946
rect 12029 5912 12035 5929
rect 12052 5912 12058 5929
rect 12029 5904 12058 5912
rect 12552 6099 12581 6104
rect 12552 6082 12558 6099
rect 12575 6082 12581 6099
rect 12552 6065 12581 6082
rect 12552 6048 12558 6065
rect 12575 6048 12581 6065
rect 12552 6031 12581 6048
rect 12552 6014 12558 6031
rect 12575 6014 12581 6031
rect 12552 5997 12581 6014
rect 12552 5980 12558 5997
rect 12575 5980 12581 5997
rect 12552 5963 12581 5980
rect 12552 5946 12558 5963
rect 12575 5946 12581 5963
rect 12552 5929 12581 5946
rect 12552 5912 12558 5929
rect 12575 5912 12581 5929
rect 12552 5904 12581 5912
rect 12596 6099 12625 6104
rect 12596 6082 12602 6099
rect 12619 6082 12625 6099
rect 12596 6065 12625 6082
rect 12596 6048 12602 6065
rect 12619 6048 12625 6065
rect 12596 6031 12625 6048
rect 12596 6014 12602 6031
rect 12619 6014 12625 6031
rect 12596 5997 12625 6014
rect 12596 5980 12602 5997
rect 12619 5980 12625 5997
rect 12596 5963 12625 5980
rect 12596 5946 12602 5963
rect 12619 5946 12625 5963
rect 12596 5929 12625 5946
rect 12596 5912 12602 5929
rect 12619 5912 12625 5929
rect 12596 5904 12625 5912
rect 12640 6099 12669 6104
rect 12640 6082 12646 6099
rect 12663 6082 12669 6099
rect 12640 6065 12669 6082
rect 12640 6048 12646 6065
rect 12663 6048 12669 6065
rect 12640 6031 12669 6048
rect 12640 6014 12646 6031
rect 12663 6014 12669 6031
rect 12640 5997 12669 6014
rect 12640 5980 12646 5997
rect 12663 5980 12669 5997
rect 12640 5963 12669 5980
rect 12640 5946 12646 5963
rect 12663 5946 12669 5963
rect 12640 5929 12669 5946
rect 12640 5912 12646 5929
rect 12663 5912 12669 5929
rect 12640 5904 12669 5912
rect 9530 5449 9559 5454
rect 9530 5432 9536 5449
rect 9553 5432 9559 5449
rect 9530 5415 9559 5432
rect 9530 5398 9536 5415
rect 9553 5398 9559 5415
rect 9530 5381 9559 5398
rect 9530 5364 9536 5381
rect 9553 5364 9559 5381
rect 9530 5347 9559 5364
rect 9530 5330 9536 5347
rect 9553 5330 9559 5347
rect 9530 5313 9559 5330
rect 9530 5296 9536 5313
rect 9553 5296 9559 5313
rect 9530 5279 9559 5296
rect 9530 5262 9536 5279
rect 9553 5262 9559 5279
rect 9530 5254 9559 5262
rect 9574 5449 9603 5454
rect 9574 5432 9580 5449
rect 9597 5432 9603 5449
rect 9574 5415 9603 5432
rect 9574 5398 9580 5415
rect 9597 5398 9603 5415
rect 9574 5381 9603 5398
rect 9574 5364 9580 5381
rect 9597 5364 9603 5381
rect 9574 5347 9603 5364
rect 9574 5330 9580 5347
rect 9597 5330 9603 5347
rect 9574 5313 9603 5330
rect 9574 5296 9580 5313
rect 9597 5296 9603 5313
rect 9574 5279 9603 5296
rect 9574 5262 9580 5279
rect 9597 5262 9603 5279
rect 9574 5254 9603 5262
rect 9618 5449 9647 5454
rect 9618 5432 9624 5449
rect 9641 5432 9647 5449
rect 9618 5415 9647 5432
rect 9618 5398 9624 5415
rect 9641 5398 9647 5415
rect 9618 5381 9647 5398
rect 9618 5364 9624 5381
rect 9641 5364 9647 5381
rect 9618 5347 9647 5364
rect 9618 5330 9624 5347
rect 9641 5330 9647 5347
rect 9618 5313 9647 5330
rect 9618 5296 9624 5313
rect 9641 5296 9647 5313
rect 9618 5279 9647 5296
rect 9618 5262 9624 5279
rect 9641 5262 9647 5279
rect 9618 5254 9647 5262
rect 10141 5449 10170 5454
rect 10141 5432 10147 5449
rect 10164 5432 10170 5449
rect 10141 5415 10170 5432
rect 10141 5398 10147 5415
rect 10164 5398 10170 5415
rect 10141 5381 10170 5398
rect 10141 5364 10147 5381
rect 10164 5364 10170 5381
rect 10141 5347 10170 5364
rect 10141 5330 10147 5347
rect 10164 5330 10170 5347
rect 10141 5313 10170 5330
rect 10141 5296 10147 5313
rect 10164 5296 10170 5313
rect 10141 5279 10170 5296
rect 10141 5262 10147 5279
rect 10164 5262 10170 5279
rect 10141 5254 10170 5262
rect 10185 5449 10214 5454
rect 10185 5432 10191 5449
rect 10208 5432 10214 5449
rect 10185 5415 10214 5432
rect 10185 5398 10191 5415
rect 10208 5398 10214 5415
rect 10185 5381 10214 5398
rect 10185 5364 10191 5381
rect 10208 5364 10214 5381
rect 10185 5347 10214 5364
rect 10185 5330 10191 5347
rect 10208 5330 10214 5347
rect 10185 5313 10214 5330
rect 10185 5296 10191 5313
rect 10208 5296 10214 5313
rect 10185 5279 10214 5296
rect 10185 5262 10191 5279
rect 10208 5262 10214 5279
rect 10185 5254 10214 5262
rect 10229 5449 10258 5454
rect 10229 5432 10235 5449
rect 10252 5432 10258 5449
rect 10229 5415 10258 5432
rect 10229 5398 10235 5415
rect 10252 5398 10258 5415
rect 10229 5381 10258 5398
rect 10229 5364 10235 5381
rect 10252 5364 10258 5381
rect 10229 5347 10258 5364
rect 10229 5330 10235 5347
rect 10252 5330 10258 5347
rect 10229 5313 10258 5330
rect 10229 5296 10235 5313
rect 10252 5296 10258 5313
rect 10229 5279 10258 5296
rect 10229 5262 10235 5279
rect 10252 5262 10258 5279
rect 10229 5254 10258 5262
rect 10752 5449 10781 5454
rect 10752 5432 10758 5449
rect 10775 5432 10781 5449
rect 10752 5415 10781 5432
rect 10752 5398 10758 5415
rect 10775 5398 10781 5415
rect 10752 5381 10781 5398
rect 10752 5364 10758 5381
rect 10775 5364 10781 5381
rect 10752 5347 10781 5364
rect 10752 5330 10758 5347
rect 10775 5330 10781 5347
rect 10752 5313 10781 5330
rect 10752 5296 10758 5313
rect 10775 5296 10781 5313
rect 10752 5279 10781 5296
rect 10752 5262 10758 5279
rect 10775 5262 10781 5279
rect 10752 5254 10781 5262
rect 10796 5449 10825 5454
rect 10796 5432 10802 5449
rect 10819 5432 10825 5449
rect 10796 5415 10825 5432
rect 10796 5398 10802 5415
rect 10819 5398 10825 5415
rect 10796 5381 10825 5398
rect 10796 5364 10802 5381
rect 10819 5364 10825 5381
rect 10796 5347 10825 5364
rect 10796 5330 10802 5347
rect 10819 5330 10825 5347
rect 10796 5313 10825 5330
rect 10796 5296 10802 5313
rect 10819 5296 10825 5313
rect 10796 5279 10825 5296
rect 10796 5262 10802 5279
rect 10819 5262 10825 5279
rect 10796 5254 10825 5262
rect 10840 5449 10869 5454
rect 10840 5432 10846 5449
rect 10863 5432 10869 5449
rect 10840 5415 10869 5432
rect 10840 5398 10846 5415
rect 10863 5398 10869 5415
rect 10840 5381 10869 5398
rect 10840 5364 10846 5381
rect 10863 5364 10869 5381
rect 10840 5347 10869 5364
rect 10840 5330 10846 5347
rect 10863 5330 10869 5347
rect 10840 5313 10869 5330
rect 10840 5296 10846 5313
rect 10863 5296 10869 5313
rect 10840 5279 10869 5296
rect 10840 5262 10846 5279
rect 10863 5262 10869 5279
rect 10840 5254 10869 5262
rect 11330 5449 11359 5454
rect 11330 5432 11336 5449
rect 11353 5432 11359 5449
rect 11330 5415 11359 5432
rect 11330 5398 11336 5415
rect 11353 5398 11359 5415
rect 11330 5381 11359 5398
rect 11330 5364 11336 5381
rect 11353 5364 11359 5381
rect 11330 5347 11359 5364
rect 11330 5330 11336 5347
rect 11353 5330 11359 5347
rect 11330 5313 11359 5330
rect 11330 5296 11336 5313
rect 11353 5296 11359 5313
rect 11330 5279 11359 5296
rect 11330 5262 11336 5279
rect 11353 5262 11359 5279
rect 11330 5254 11359 5262
rect 11374 5449 11403 5454
rect 11374 5432 11380 5449
rect 11397 5432 11403 5449
rect 11374 5415 11403 5432
rect 11374 5398 11380 5415
rect 11397 5398 11403 5415
rect 11374 5381 11403 5398
rect 11374 5364 11380 5381
rect 11397 5364 11403 5381
rect 11374 5347 11403 5364
rect 11374 5330 11380 5347
rect 11397 5330 11403 5347
rect 11374 5313 11403 5330
rect 11374 5296 11380 5313
rect 11397 5296 11403 5313
rect 11374 5279 11403 5296
rect 11374 5262 11380 5279
rect 11397 5262 11403 5279
rect 11374 5254 11403 5262
rect 11418 5449 11447 5454
rect 11418 5432 11424 5449
rect 11441 5432 11447 5449
rect 11418 5415 11447 5432
rect 11418 5398 11424 5415
rect 11441 5398 11447 5415
rect 11418 5381 11447 5398
rect 11418 5364 11424 5381
rect 11441 5364 11447 5381
rect 11418 5347 11447 5364
rect 11418 5330 11424 5347
rect 11441 5330 11447 5347
rect 11418 5313 11447 5330
rect 11418 5296 11424 5313
rect 11441 5296 11447 5313
rect 11418 5279 11447 5296
rect 11418 5262 11424 5279
rect 11441 5262 11447 5279
rect 11418 5254 11447 5262
rect 11941 5449 11970 5454
rect 11941 5432 11947 5449
rect 11964 5432 11970 5449
rect 11941 5415 11970 5432
rect 11941 5398 11947 5415
rect 11964 5398 11970 5415
rect 11941 5381 11970 5398
rect 11941 5364 11947 5381
rect 11964 5364 11970 5381
rect 11941 5347 11970 5364
rect 11941 5330 11947 5347
rect 11964 5330 11970 5347
rect 11941 5313 11970 5330
rect 11941 5296 11947 5313
rect 11964 5296 11970 5313
rect 11941 5279 11970 5296
rect 11941 5262 11947 5279
rect 11964 5262 11970 5279
rect 11941 5254 11970 5262
rect 11985 5449 12014 5454
rect 11985 5432 11991 5449
rect 12008 5432 12014 5449
rect 11985 5415 12014 5432
rect 11985 5398 11991 5415
rect 12008 5398 12014 5415
rect 11985 5381 12014 5398
rect 11985 5364 11991 5381
rect 12008 5364 12014 5381
rect 11985 5347 12014 5364
rect 11985 5330 11991 5347
rect 12008 5330 12014 5347
rect 11985 5313 12014 5330
rect 11985 5296 11991 5313
rect 12008 5296 12014 5313
rect 11985 5279 12014 5296
rect 11985 5262 11991 5279
rect 12008 5262 12014 5279
rect 11985 5254 12014 5262
rect 12029 5449 12058 5454
rect 12029 5432 12035 5449
rect 12052 5432 12058 5449
rect 12029 5415 12058 5432
rect 12029 5398 12035 5415
rect 12052 5398 12058 5415
rect 12029 5381 12058 5398
rect 12029 5364 12035 5381
rect 12052 5364 12058 5381
rect 12029 5347 12058 5364
rect 12029 5330 12035 5347
rect 12052 5330 12058 5347
rect 12029 5313 12058 5330
rect 12029 5296 12035 5313
rect 12052 5296 12058 5313
rect 12029 5279 12058 5296
rect 12029 5262 12035 5279
rect 12052 5262 12058 5279
rect 12029 5254 12058 5262
rect 12552 5449 12581 5454
rect 12552 5432 12558 5449
rect 12575 5432 12581 5449
rect 12552 5415 12581 5432
rect 12552 5398 12558 5415
rect 12575 5398 12581 5415
rect 12552 5381 12581 5398
rect 12552 5364 12558 5381
rect 12575 5364 12581 5381
rect 12552 5347 12581 5364
rect 12552 5330 12558 5347
rect 12575 5330 12581 5347
rect 12552 5313 12581 5330
rect 12552 5296 12558 5313
rect 12575 5296 12581 5313
rect 12552 5279 12581 5296
rect 12552 5262 12558 5279
rect 12575 5262 12581 5279
rect 12552 5254 12581 5262
rect 12596 5449 12625 5454
rect 12596 5432 12602 5449
rect 12619 5432 12625 5449
rect 12596 5415 12625 5432
rect 12596 5398 12602 5415
rect 12619 5398 12625 5415
rect 12596 5381 12625 5398
rect 12596 5364 12602 5381
rect 12619 5364 12625 5381
rect 12596 5347 12625 5364
rect 12596 5330 12602 5347
rect 12619 5330 12625 5347
rect 12596 5313 12625 5330
rect 12596 5296 12602 5313
rect 12619 5296 12625 5313
rect 12596 5279 12625 5296
rect 12596 5262 12602 5279
rect 12619 5262 12625 5279
rect 12596 5254 12625 5262
rect 12640 5449 12669 5454
rect 12640 5432 12646 5449
rect 12663 5432 12669 5449
rect 12640 5415 12669 5432
rect 12640 5398 12646 5415
rect 12663 5398 12669 5415
rect 12640 5381 12669 5398
rect 12640 5364 12646 5381
rect 12663 5364 12669 5381
rect 12640 5347 12669 5364
rect 12640 5330 12646 5347
rect 12663 5330 12669 5347
rect 12640 5313 12669 5330
rect 12640 5296 12646 5313
rect 12663 5296 12669 5313
rect 12640 5279 12669 5296
rect 12640 5262 12646 5279
rect 12663 5262 12669 5279
rect 12640 5254 12669 5262
rect 9530 4809 9559 4814
rect 9530 4792 9536 4809
rect 9553 4792 9559 4809
rect 9530 4775 9559 4792
rect 9530 4758 9536 4775
rect 9553 4758 9559 4775
rect 9530 4741 9559 4758
rect 9530 4724 9536 4741
rect 9553 4724 9559 4741
rect 9530 4707 9559 4724
rect 9530 4690 9536 4707
rect 9553 4690 9559 4707
rect 9530 4673 9559 4690
rect 9530 4656 9536 4673
rect 9553 4656 9559 4673
rect 9530 4639 9559 4656
rect 9530 4622 9536 4639
rect 9553 4622 9559 4639
rect 9530 4614 9559 4622
rect 9574 4809 9603 4814
rect 9574 4792 9580 4809
rect 9597 4792 9603 4809
rect 9574 4775 9603 4792
rect 9574 4758 9580 4775
rect 9597 4758 9603 4775
rect 9574 4741 9603 4758
rect 9574 4724 9580 4741
rect 9597 4724 9603 4741
rect 9574 4707 9603 4724
rect 9574 4690 9580 4707
rect 9597 4690 9603 4707
rect 9574 4673 9603 4690
rect 9574 4656 9580 4673
rect 9597 4656 9603 4673
rect 9574 4639 9603 4656
rect 9574 4622 9580 4639
rect 9597 4622 9603 4639
rect 9574 4614 9603 4622
rect 9618 4809 9647 4814
rect 9618 4792 9624 4809
rect 9641 4792 9647 4809
rect 9618 4775 9647 4792
rect 9618 4758 9624 4775
rect 9641 4758 9647 4775
rect 9618 4741 9647 4758
rect 9618 4724 9624 4741
rect 9641 4724 9647 4741
rect 9618 4707 9647 4724
rect 9618 4690 9624 4707
rect 9641 4690 9647 4707
rect 9618 4673 9647 4690
rect 9618 4656 9624 4673
rect 9641 4656 9647 4673
rect 9618 4639 9647 4656
rect 9618 4622 9624 4639
rect 9641 4622 9647 4639
rect 9618 4614 9647 4622
rect 10141 4809 10170 4814
rect 10141 4792 10147 4809
rect 10164 4792 10170 4809
rect 10141 4775 10170 4792
rect 10141 4758 10147 4775
rect 10164 4758 10170 4775
rect 10141 4741 10170 4758
rect 10141 4724 10147 4741
rect 10164 4724 10170 4741
rect 10141 4707 10170 4724
rect 10141 4690 10147 4707
rect 10164 4690 10170 4707
rect 10141 4673 10170 4690
rect 10141 4656 10147 4673
rect 10164 4656 10170 4673
rect 10141 4639 10170 4656
rect 10141 4622 10147 4639
rect 10164 4622 10170 4639
rect 10141 4614 10170 4622
rect 10185 4809 10214 4814
rect 10185 4792 10191 4809
rect 10208 4792 10214 4809
rect 10185 4775 10214 4792
rect 10185 4758 10191 4775
rect 10208 4758 10214 4775
rect 10185 4741 10214 4758
rect 10185 4724 10191 4741
rect 10208 4724 10214 4741
rect 10185 4707 10214 4724
rect 10185 4690 10191 4707
rect 10208 4690 10214 4707
rect 10185 4673 10214 4690
rect 10185 4656 10191 4673
rect 10208 4656 10214 4673
rect 10185 4639 10214 4656
rect 10185 4622 10191 4639
rect 10208 4622 10214 4639
rect 10185 4614 10214 4622
rect 10229 4809 10258 4814
rect 10229 4792 10235 4809
rect 10252 4792 10258 4809
rect 10229 4775 10258 4792
rect 10229 4758 10235 4775
rect 10252 4758 10258 4775
rect 10229 4741 10258 4758
rect 10229 4724 10235 4741
rect 10252 4724 10258 4741
rect 10229 4707 10258 4724
rect 10229 4690 10235 4707
rect 10252 4690 10258 4707
rect 10229 4673 10258 4690
rect 10229 4656 10235 4673
rect 10252 4656 10258 4673
rect 10229 4639 10258 4656
rect 10229 4622 10235 4639
rect 10252 4622 10258 4639
rect 10229 4614 10258 4622
rect 10752 4809 10781 4814
rect 10752 4792 10758 4809
rect 10775 4792 10781 4809
rect 10752 4775 10781 4792
rect 10752 4758 10758 4775
rect 10775 4758 10781 4775
rect 10752 4741 10781 4758
rect 10752 4724 10758 4741
rect 10775 4724 10781 4741
rect 10752 4707 10781 4724
rect 10752 4690 10758 4707
rect 10775 4690 10781 4707
rect 10752 4673 10781 4690
rect 10752 4656 10758 4673
rect 10775 4656 10781 4673
rect 10752 4639 10781 4656
rect 10752 4622 10758 4639
rect 10775 4622 10781 4639
rect 10752 4614 10781 4622
rect 10796 4809 10825 4814
rect 10796 4792 10802 4809
rect 10819 4792 10825 4809
rect 10796 4775 10825 4792
rect 10796 4758 10802 4775
rect 10819 4758 10825 4775
rect 10796 4741 10825 4758
rect 10796 4724 10802 4741
rect 10819 4724 10825 4741
rect 10796 4707 10825 4724
rect 10796 4690 10802 4707
rect 10819 4690 10825 4707
rect 10796 4673 10825 4690
rect 10796 4656 10802 4673
rect 10819 4656 10825 4673
rect 10796 4639 10825 4656
rect 10796 4622 10802 4639
rect 10819 4622 10825 4639
rect 10796 4614 10825 4622
rect 10840 4809 10869 4814
rect 10840 4792 10846 4809
rect 10863 4792 10869 4809
rect 10840 4775 10869 4792
rect 10840 4758 10846 4775
rect 10863 4758 10869 4775
rect 10840 4741 10869 4758
rect 10840 4724 10846 4741
rect 10863 4724 10869 4741
rect 10840 4707 10869 4724
rect 10840 4690 10846 4707
rect 10863 4690 10869 4707
rect 10840 4673 10869 4690
rect 10840 4656 10846 4673
rect 10863 4656 10869 4673
rect 10840 4639 10869 4656
rect 10840 4622 10846 4639
rect 10863 4622 10869 4639
rect 10840 4614 10869 4622
rect 11330 4809 11359 4814
rect 11330 4792 11336 4809
rect 11353 4792 11359 4809
rect 11330 4775 11359 4792
rect 11330 4758 11336 4775
rect 11353 4758 11359 4775
rect 11330 4741 11359 4758
rect 11330 4724 11336 4741
rect 11353 4724 11359 4741
rect 11330 4707 11359 4724
rect 11330 4690 11336 4707
rect 11353 4690 11359 4707
rect 11330 4673 11359 4690
rect 11330 4656 11336 4673
rect 11353 4656 11359 4673
rect 11330 4639 11359 4656
rect 11330 4622 11336 4639
rect 11353 4622 11359 4639
rect 11330 4614 11359 4622
rect 11374 4809 11403 4814
rect 11374 4792 11380 4809
rect 11397 4792 11403 4809
rect 11374 4775 11403 4792
rect 11374 4758 11380 4775
rect 11397 4758 11403 4775
rect 11374 4741 11403 4758
rect 11374 4724 11380 4741
rect 11397 4724 11403 4741
rect 11374 4707 11403 4724
rect 11374 4690 11380 4707
rect 11397 4690 11403 4707
rect 11374 4673 11403 4690
rect 11374 4656 11380 4673
rect 11397 4656 11403 4673
rect 11374 4639 11403 4656
rect 11374 4622 11380 4639
rect 11397 4622 11403 4639
rect 11374 4614 11403 4622
rect 11418 4809 11447 4814
rect 11418 4792 11424 4809
rect 11441 4792 11447 4809
rect 11418 4775 11447 4792
rect 11418 4758 11424 4775
rect 11441 4758 11447 4775
rect 11418 4741 11447 4758
rect 11418 4724 11424 4741
rect 11441 4724 11447 4741
rect 11418 4707 11447 4724
rect 11418 4690 11424 4707
rect 11441 4690 11447 4707
rect 11418 4673 11447 4690
rect 11418 4656 11424 4673
rect 11441 4656 11447 4673
rect 11418 4639 11447 4656
rect 11418 4622 11424 4639
rect 11441 4622 11447 4639
rect 11418 4614 11447 4622
rect 11941 4809 11970 4814
rect 11941 4792 11947 4809
rect 11964 4792 11970 4809
rect 11941 4775 11970 4792
rect 11941 4758 11947 4775
rect 11964 4758 11970 4775
rect 11941 4741 11970 4758
rect 11941 4724 11947 4741
rect 11964 4724 11970 4741
rect 11941 4707 11970 4724
rect 11941 4690 11947 4707
rect 11964 4690 11970 4707
rect 11941 4673 11970 4690
rect 11941 4656 11947 4673
rect 11964 4656 11970 4673
rect 11941 4639 11970 4656
rect 11941 4622 11947 4639
rect 11964 4622 11970 4639
rect 11941 4614 11970 4622
rect 11985 4809 12014 4814
rect 11985 4792 11991 4809
rect 12008 4792 12014 4809
rect 11985 4775 12014 4792
rect 11985 4758 11991 4775
rect 12008 4758 12014 4775
rect 11985 4741 12014 4758
rect 11985 4724 11991 4741
rect 12008 4724 12014 4741
rect 11985 4707 12014 4724
rect 11985 4690 11991 4707
rect 12008 4690 12014 4707
rect 11985 4673 12014 4690
rect 11985 4656 11991 4673
rect 12008 4656 12014 4673
rect 11985 4639 12014 4656
rect 11985 4622 11991 4639
rect 12008 4622 12014 4639
rect 11985 4614 12014 4622
rect 12029 4809 12058 4814
rect 12029 4792 12035 4809
rect 12052 4792 12058 4809
rect 12029 4775 12058 4792
rect 12029 4758 12035 4775
rect 12052 4758 12058 4775
rect 12029 4741 12058 4758
rect 12029 4724 12035 4741
rect 12052 4724 12058 4741
rect 12029 4707 12058 4724
rect 12029 4690 12035 4707
rect 12052 4690 12058 4707
rect 12029 4673 12058 4690
rect 12029 4656 12035 4673
rect 12052 4656 12058 4673
rect 12029 4639 12058 4656
rect 12029 4622 12035 4639
rect 12052 4622 12058 4639
rect 12029 4614 12058 4622
rect 12552 4809 12581 4814
rect 12552 4792 12558 4809
rect 12575 4792 12581 4809
rect 12552 4775 12581 4792
rect 12552 4758 12558 4775
rect 12575 4758 12581 4775
rect 12552 4741 12581 4758
rect 12552 4724 12558 4741
rect 12575 4724 12581 4741
rect 12552 4707 12581 4724
rect 12552 4690 12558 4707
rect 12575 4690 12581 4707
rect 12552 4673 12581 4690
rect 12552 4656 12558 4673
rect 12575 4656 12581 4673
rect 12552 4639 12581 4656
rect 12552 4622 12558 4639
rect 12575 4622 12581 4639
rect 12552 4614 12581 4622
rect 12596 4809 12625 4814
rect 12596 4792 12602 4809
rect 12619 4792 12625 4809
rect 12596 4775 12625 4792
rect 12596 4758 12602 4775
rect 12619 4758 12625 4775
rect 12596 4741 12625 4758
rect 12596 4724 12602 4741
rect 12619 4724 12625 4741
rect 12596 4707 12625 4724
rect 12596 4690 12602 4707
rect 12619 4690 12625 4707
rect 12596 4673 12625 4690
rect 12596 4656 12602 4673
rect 12619 4656 12625 4673
rect 12596 4639 12625 4656
rect 12596 4622 12602 4639
rect 12619 4622 12625 4639
rect 12596 4614 12625 4622
rect 12640 4809 12669 4814
rect 12640 4792 12646 4809
rect 12663 4792 12669 4809
rect 12640 4775 12669 4792
rect 12640 4758 12646 4775
rect 12663 4758 12669 4775
rect 12640 4741 12669 4758
rect 12640 4724 12646 4741
rect 12663 4724 12669 4741
rect 12640 4707 12669 4724
rect 12640 4690 12646 4707
rect 12663 4690 12669 4707
rect 12640 4673 12669 4690
rect 12640 4656 12646 4673
rect 12663 4656 12669 4673
rect 12640 4639 12669 4656
rect 12640 4622 12646 4639
rect 12663 4622 12669 4639
rect 12640 4614 12669 4622
<< ndiffc >>
rect 10067 7646 10084 7663
rect 10067 7612 10084 7629
rect 10067 7578 10084 7595
rect 10147 7646 10164 7663
rect 10147 7612 10164 7629
rect 10147 7578 10164 7595
rect 10191 7646 10208 7663
rect 10191 7612 10208 7629
rect 10191 7578 10208 7595
rect 10235 7646 10252 7663
rect 10235 7612 10252 7629
rect 10235 7578 10252 7595
rect 10315 7646 10332 7663
rect 10315 7612 10332 7629
rect 10315 7578 10332 7595
rect 10678 7646 10695 7663
rect 10678 7612 10695 7629
rect 10678 7578 10695 7595
rect 10758 7646 10775 7663
rect 10758 7612 10775 7629
rect 10758 7578 10775 7595
rect 10802 7646 10819 7663
rect 10802 7612 10819 7629
rect 10802 7578 10819 7595
rect 10846 7646 10863 7663
rect 10846 7612 10863 7629
rect 10846 7578 10863 7595
rect 10926 7646 10943 7663
rect 10926 7612 10943 7629
rect 10926 7578 10943 7595
rect 11256 7646 11273 7663
rect 11256 7612 11273 7629
rect 11256 7578 11273 7595
rect 11336 7646 11353 7663
rect 11336 7612 11353 7629
rect 11336 7578 11353 7595
rect 11380 7646 11397 7663
rect 11380 7612 11397 7629
rect 11380 7578 11397 7595
rect 11424 7646 11441 7663
rect 11424 7612 11441 7629
rect 11424 7578 11441 7595
rect 11504 7646 11521 7663
rect 11504 7612 11521 7629
rect 11504 7578 11521 7595
rect 11867 7646 11884 7663
rect 11867 7612 11884 7629
rect 11867 7578 11884 7595
rect 11947 7646 11964 7663
rect 11947 7612 11964 7629
rect 11947 7578 11964 7595
rect 11991 7646 12008 7663
rect 11991 7612 12008 7629
rect 11991 7578 12008 7595
rect 12035 7646 12052 7663
rect 12035 7612 12052 7629
rect 12035 7578 12052 7595
rect 12115 7646 12132 7663
rect 12115 7612 12132 7629
rect 12115 7578 12132 7595
rect 12478 7646 12495 7663
rect 12478 7612 12495 7629
rect 12478 7578 12495 7595
rect 12558 7646 12575 7663
rect 12558 7612 12575 7629
rect 12558 7578 12575 7595
rect 12602 7646 12619 7663
rect 12602 7612 12619 7629
rect 12602 7578 12619 7595
rect 12646 7646 12663 7663
rect 12646 7612 12663 7629
rect 12646 7578 12663 7595
rect 12726 7646 12743 7663
rect 12726 7612 12743 7629
rect 12726 7578 12743 7595
rect 9456 6996 9473 7013
rect 9456 6962 9473 6979
rect 9456 6928 9473 6945
rect 9536 6996 9553 7013
rect 9536 6962 9553 6979
rect 9536 6928 9553 6945
rect 9580 6996 9597 7013
rect 9580 6962 9597 6979
rect 9580 6928 9597 6945
rect 9624 6996 9641 7013
rect 9624 6962 9641 6979
rect 9624 6928 9641 6945
rect 9704 6996 9721 7013
rect 9704 6962 9721 6979
rect 9704 6928 9721 6945
rect 10067 6996 10084 7013
rect 10067 6962 10084 6979
rect 10067 6928 10084 6945
rect 10147 6996 10164 7013
rect 10147 6962 10164 6979
rect 10147 6928 10164 6945
rect 10191 6996 10208 7013
rect 10191 6962 10208 6979
rect 10191 6928 10208 6945
rect 10235 6996 10252 7013
rect 10235 6962 10252 6979
rect 10235 6928 10252 6945
rect 10315 6996 10332 7013
rect 10315 6962 10332 6979
rect 10315 6928 10332 6945
rect 10678 6996 10695 7013
rect 10678 6962 10695 6979
rect 10678 6928 10695 6945
rect 10758 6996 10775 7013
rect 10758 6962 10775 6979
rect 10758 6928 10775 6945
rect 10802 6996 10819 7013
rect 10802 6962 10819 6979
rect 10802 6928 10819 6945
rect 10846 6996 10863 7013
rect 10846 6962 10863 6979
rect 10846 6928 10863 6945
rect 10926 6996 10943 7013
rect 10926 6962 10943 6979
rect 10926 6928 10943 6945
rect 11256 6996 11273 7013
rect 11256 6962 11273 6979
rect 11256 6928 11273 6945
rect 11336 6996 11353 7013
rect 11336 6962 11353 6979
rect 11336 6928 11353 6945
rect 11380 6996 11397 7013
rect 11380 6962 11397 6979
rect 11380 6928 11397 6945
rect 11424 6996 11441 7013
rect 11424 6962 11441 6979
rect 11424 6928 11441 6945
rect 11504 6996 11521 7013
rect 11504 6962 11521 6979
rect 11504 6928 11521 6945
rect 11867 6996 11884 7013
rect 11867 6962 11884 6979
rect 11867 6928 11884 6945
rect 11947 6996 11964 7013
rect 11947 6962 11964 6979
rect 11947 6928 11964 6945
rect 11991 6996 12008 7013
rect 11991 6962 12008 6979
rect 11991 6928 12008 6945
rect 12035 6996 12052 7013
rect 12035 6962 12052 6979
rect 12035 6928 12052 6945
rect 12115 6996 12132 7013
rect 12115 6962 12132 6979
rect 12115 6928 12132 6945
rect 12478 6996 12495 7013
rect 12478 6962 12495 6979
rect 12478 6928 12495 6945
rect 12558 6996 12575 7013
rect 12558 6962 12575 6979
rect 12558 6928 12575 6945
rect 12602 6996 12619 7013
rect 12602 6962 12619 6979
rect 12602 6928 12619 6945
rect 12646 6996 12663 7013
rect 12646 6962 12663 6979
rect 12646 6928 12663 6945
rect 12726 6996 12743 7013
rect 12726 6962 12743 6979
rect 12726 6928 12743 6945
rect 9456 6356 9473 6373
rect 9456 6322 9473 6339
rect 9456 6288 9473 6305
rect 9536 6356 9553 6373
rect 9536 6322 9553 6339
rect 9536 6288 9553 6305
rect 9580 6356 9597 6373
rect 9580 6322 9597 6339
rect 9580 6288 9597 6305
rect 9624 6356 9641 6373
rect 9624 6322 9641 6339
rect 9624 6288 9641 6305
rect 9704 6356 9721 6373
rect 9704 6322 9721 6339
rect 9704 6288 9721 6305
rect 10067 6356 10084 6373
rect 10067 6322 10084 6339
rect 10067 6288 10084 6305
rect 10147 6356 10164 6373
rect 10147 6322 10164 6339
rect 10147 6288 10164 6305
rect 10191 6356 10208 6373
rect 10191 6322 10208 6339
rect 10191 6288 10208 6305
rect 10235 6356 10252 6373
rect 10235 6322 10252 6339
rect 10235 6288 10252 6305
rect 10315 6356 10332 6373
rect 10315 6322 10332 6339
rect 10315 6288 10332 6305
rect 10678 6356 10695 6373
rect 10678 6322 10695 6339
rect 10678 6288 10695 6305
rect 10758 6356 10775 6373
rect 10758 6322 10775 6339
rect 10758 6288 10775 6305
rect 10802 6356 10819 6373
rect 10802 6322 10819 6339
rect 10802 6288 10819 6305
rect 10846 6356 10863 6373
rect 10846 6322 10863 6339
rect 10846 6288 10863 6305
rect 10926 6356 10943 6373
rect 10926 6322 10943 6339
rect 10926 6288 10943 6305
rect 11256 6356 11273 6373
rect 11256 6322 11273 6339
rect 11256 6288 11273 6305
rect 11336 6356 11353 6373
rect 11336 6322 11353 6339
rect 11336 6288 11353 6305
rect 11380 6356 11397 6373
rect 11380 6322 11397 6339
rect 11380 6288 11397 6305
rect 11424 6356 11441 6373
rect 11424 6322 11441 6339
rect 11424 6288 11441 6305
rect 11504 6356 11521 6373
rect 11504 6322 11521 6339
rect 11504 6288 11521 6305
rect 11867 6356 11884 6373
rect 11867 6322 11884 6339
rect 11867 6288 11884 6305
rect 11947 6356 11964 6373
rect 11947 6322 11964 6339
rect 11947 6288 11964 6305
rect 11991 6356 12008 6373
rect 11991 6322 12008 6339
rect 11991 6288 12008 6305
rect 12035 6356 12052 6373
rect 12035 6322 12052 6339
rect 12035 6288 12052 6305
rect 12115 6356 12132 6373
rect 12115 6322 12132 6339
rect 12115 6288 12132 6305
rect 12478 6356 12495 6373
rect 12478 6322 12495 6339
rect 12478 6288 12495 6305
rect 12558 6356 12575 6373
rect 12558 6322 12575 6339
rect 12558 6288 12575 6305
rect 12602 6356 12619 6373
rect 12602 6322 12619 6339
rect 12602 6288 12619 6305
rect 12646 6356 12663 6373
rect 12646 6322 12663 6339
rect 12646 6288 12663 6305
rect 12726 6356 12743 6373
rect 12726 6322 12743 6339
rect 12726 6288 12743 6305
rect 9456 5706 9473 5723
rect 9456 5672 9473 5689
rect 9456 5638 9473 5655
rect 9536 5706 9553 5723
rect 9536 5672 9553 5689
rect 9536 5638 9553 5655
rect 9580 5706 9597 5723
rect 9580 5672 9597 5689
rect 9580 5638 9597 5655
rect 9624 5706 9641 5723
rect 9624 5672 9641 5689
rect 9624 5638 9641 5655
rect 9704 5706 9721 5723
rect 9704 5672 9721 5689
rect 9704 5638 9721 5655
rect 10067 5706 10084 5723
rect 10067 5672 10084 5689
rect 10067 5638 10084 5655
rect 10147 5706 10164 5723
rect 10147 5672 10164 5689
rect 10147 5638 10164 5655
rect 10191 5706 10208 5723
rect 10191 5672 10208 5689
rect 10191 5638 10208 5655
rect 10235 5706 10252 5723
rect 10235 5672 10252 5689
rect 10235 5638 10252 5655
rect 10315 5706 10332 5723
rect 10315 5672 10332 5689
rect 10315 5638 10332 5655
rect 10678 5706 10695 5723
rect 10678 5672 10695 5689
rect 10678 5638 10695 5655
rect 10758 5706 10775 5723
rect 10758 5672 10775 5689
rect 10758 5638 10775 5655
rect 10802 5706 10819 5723
rect 10802 5672 10819 5689
rect 10802 5638 10819 5655
rect 10846 5706 10863 5723
rect 10846 5672 10863 5689
rect 10846 5638 10863 5655
rect 10926 5706 10943 5723
rect 10926 5672 10943 5689
rect 10926 5638 10943 5655
rect 11256 5706 11273 5723
rect 11256 5672 11273 5689
rect 11256 5638 11273 5655
rect 11336 5706 11353 5723
rect 11336 5672 11353 5689
rect 11336 5638 11353 5655
rect 11380 5706 11397 5723
rect 11380 5672 11397 5689
rect 11380 5638 11397 5655
rect 11424 5706 11441 5723
rect 11424 5672 11441 5689
rect 11424 5638 11441 5655
rect 11504 5706 11521 5723
rect 11504 5672 11521 5689
rect 11504 5638 11521 5655
rect 11867 5706 11884 5723
rect 11867 5672 11884 5689
rect 11867 5638 11884 5655
rect 11947 5706 11964 5723
rect 11947 5672 11964 5689
rect 11947 5638 11964 5655
rect 11991 5706 12008 5723
rect 11991 5672 12008 5689
rect 11991 5638 12008 5655
rect 12035 5706 12052 5723
rect 12035 5672 12052 5689
rect 12035 5638 12052 5655
rect 12115 5706 12132 5723
rect 12115 5672 12132 5689
rect 12115 5638 12132 5655
rect 12478 5706 12495 5723
rect 12478 5672 12495 5689
rect 12478 5638 12495 5655
rect 12558 5706 12575 5723
rect 12558 5672 12575 5689
rect 12558 5638 12575 5655
rect 12602 5706 12619 5723
rect 12602 5672 12619 5689
rect 12602 5638 12619 5655
rect 12646 5706 12663 5723
rect 12646 5672 12663 5689
rect 12646 5638 12663 5655
rect 12726 5706 12743 5723
rect 12726 5672 12743 5689
rect 12726 5638 12743 5655
rect 9456 5056 9473 5073
rect 9456 5022 9473 5039
rect 9456 4988 9473 5005
rect 9536 5056 9553 5073
rect 9536 5022 9553 5039
rect 9536 4988 9553 5005
rect 9580 5056 9597 5073
rect 9580 5022 9597 5039
rect 9580 4988 9597 5005
rect 9624 5056 9641 5073
rect 9624 5022 9641 5039
rect 9624 4988 9641 5005
rect 9704 5056 9721 5073
rect 9704 5022 9721 5039
rect 9704 4988 9721 5005
rect 10067 5056 10084 5073
rect 10067 5022 10084 5039
rect 10067 4988 10084 5005
rect 10147 5056 10164 5073
rect 10147 5022 10164 5039
rect 10147 4988 10164 5005
rect 10191 5056 10208 5073
rect 10191 5022 10208 5039
rect 10191 4988 10208 5005
rect 10235 5056 10252 5073
rect 10235 5022 10252 5039
rect 10235 4988 10252 5005
rect 10315 5056 10332 5073
rect 10315 5022 10332 5039
rect 10315 4988 10332 5005
rect 10678 5056 10695 5073
rect 10678 5022 10695 5039
rect 10678 4988 10695 5005
rect 10758 5056 10775 5073
rect 10758 5022 10775 5039
rect 10758 4988 10775 5005
rect 10802 5056 10819 5073
rect 10802 5022 10819 5039
rect 10802 4988 10819 5005
rect 10846 5056 10863 5073
rect 10846 5022 10863 5039
rect 10846 4988 10863 5005
rect 10926 5056 10943 5073
rect 10926 5022 10943 5039
rect 10926 4988 10943 5005
rect 11256 5056 11273 5073
rect 11256 5022 11273 5039
rect 11256 4988 11273 5005
rect 11336 5056 11353 5073
rect 11336 5022 11353 5039
rect 11336 4988 11353 5005
rect 11380 5056 11397 5073
rect 11380 5022 11397 5039
rect 11380 4988 11397 5005
rect 11424 5056 11441 5073
rect 11424 5022 11441 5039
rect 11424 4988 11441 5005
rect 11504 5056 11521 5073
rect 11504 5022 11521 5039
rect 11504 4988 11521 5005
rect 11867 5056 11884 5073
rect 11867 5022 11884 5039
rect 11867 4988 11884 5005
rect 11947 5056 11964 5073
rect 11947 5022 11964 5039
rect 11947 4988 11964 5005
rect 11991 5056 12008 5073
rect 11991 5022 12008 5039
rect 11991 4988 12008 5005
rect 12035 5056 12052 5073
rect 12035 5022 12052 5039
rect 12035 4988 12052 5005
rect 12115 5056 12132 5073
rect 12115 5022 12132 5039
rect 12115 4988 12132 5005
rect 12478 5056 12495 5073
rect 12478 5022 12495 5039
rect 12478 4988 12495 5005
rect 12558 5056 12575 5073
rect 12558 5022 12575 5039
rect 12558 4988 12575 5005
rect 12602 5056 12619 5073
rect 12602 5022 12619 5039
rect 12602 4988 12619 5005
rect 12646 5056 12663 5073
rect 12646 5022 12663 5039
rect 12646 4988 12663 5005
rect 12726 5056 12743 5073
rect 12726 5022 12743 5039
rect 12726 4988 12743 5005
rect 9456 4416 9473 4433
rect 9456 4382 9473 4399
rect 9456 4348 9473 4365
rect 9536 4416 9553 4433
rect 9536 4382 9553 4399
rect 9536 4348 9553 4365
rect 9580 4416 9597 4433
rect 9580 4382 9597 4399
rect 9580 4348 9597 4365
rect 9624 4416 9641 4433
rect 9624 4382 9641 4399
rect 9624 4348 9641 4365
rect 9704 4416 9721 4433
rect 9704 4382 9721 4399
rect 9704 4348 9721 4365
rect 10067 4416 10084 4433
rect 10067 4382 10084 4399
rect 10067 4348 10084 4365
rect 10147 4416 10164 4433
rect 10147 4382 10164 4399
rect 10147 4348 10164 4365
rect 10191 4416 10208 4433
rect 10191 4382 10208 4399
rect 10191 4348 10208 4365
rect 10235 4416 10252 4433
rect 10235 4382 10252 4399
rect 10235 4348 10252 4365
rect 10315 4416 10332 4433
rect 10315 4382 10332 4399
rect 10315 4348 10332 4365
rect 10678 4416 10695 4433
rect 10678 4382 10695 4399
rect 10678 4348 10695 4365
rect 10758 4416 10775 4433
rect 10758 4382 10775 4399
rect 10758 4348 10775 4365
rect 10802 4416 10819 4433
rect 10802 4382 10819 4399
rect 10802 4348 10819 4365
rect 10846 4416 10863 4433
rect 10846 4382 10863 4399
rect 10846 4348 10863 4365
rect 10926 4416 10943 4433
rect 10926 4382 10943 4399
rect 10926 4348 10943 4365
rect 11256 4416 11273 4433
rect 11256 4382 11273 4399
rect 11256 4348 11273 4365
rect 11336 4416 11353 4433
rect 11336 4382 11353 4399
rect 11336 4348 11353 4365
rect 11380 4416 11397 4433
rect 11380 4382 11397 4399
rect 11380 4348 11397 4365
rect 11424 4416 11441 4433
rect 11424 4382 11441 4399
rect 11424 4348 11441 4365
rect 11504 4416 11521 4433
rect 11504 4382 11521 4399
rect 11504 4348 11521 4365
rect 11867 4416 11884 4433
rect 11867 4382 11884 4399
rect 11867 4348 11884 4365
rect 11947 4416 11964 4433
rect 11947 4382 11964 4399
rect 11947 4348 11964 4365
rect 11991 4416 12008 4433
rect 11991 4382 12008 4399
rect 11991 4348 12008 4365
rect 12035 4416 12052 4433
rect 12035 4382 12052 4399
rect 12035 4348 12052 4365
rect 12115 4416 12132 4433
rect 12115 4382 12132 4399
rect 12115 4348 12132 4365
rect 12478 4416 12495 4433
rect 12478 4382 12495 4399
rect 12478 4348 12495 4365
rect 12558 4416 12575 4433
rect 12558 4382 12575 4399
rect 12558 4348 12575 4365
rect 12602 4416 12619 4433
rect 12602 4382 12619 4399
rect 12602 4348 12619 4365
rect 12646 4416 12663 4433
rect 12646 4382 12663 4399
rect 12646 4348 12663 4365
rect 12726 4416 12743 4433
rect 12726 4382 12743 4399
rect 12726 4348 12743 4365
<< pdiffc >>
rect 10147 8022 10164 8039
rect 10147 7988 10164 8005
rect 10147 7954 10164 7971
rect 10147 7920 10164 7937
rect 10147 7886 10164 7903
rect 10147 7852 10164 7869
rect 10191 8022 10208 8039
rect 10191 7988 10208 8005
rect 10191 7954 10208 7971
rect 10191 7920 10208 7937
rect 10191 7886 10208 7903
rect 10191 7852 10208 7869
rect 10235 8022 10252 8039
rect 10235 7988 10252 8005
rect 10235 7954 10252 7971
rect 10235 7920 10252 7937
rect 10235 7886 10252 7903
rect 10235 7852 10252 7869
rect 10758 8022 10775 8039
rect 10758 7988 10775 8005
rect 10758 7954 10775 7971
rect 10758 7920 10775 7937
rect 10758 7886 10775 7903
rect 10758 7852 10775 7869
rect 10802 8022 10819 8039
rect 10802 7988 10819 8005
rect 10802 7954 10819 7971
rect 10802 7920 10819 7937
rect 10802 7886 10819 7903
rect 10802 7852 10819 7869
rect 10846 8022 10863 8039
rect 10846 7988 10863 8005
rect 10846 7954 10863 7971
rect 10846 7920 10863 7937
rect 10846 7886 10863 7903
rect 10846 7852 10863 7869
rect 11336 8022 11353 8039
rect 11336 7988 11353 8005
rect 11336 7954 11353 7971
rect 11336 7920 11353 7937
rect 11336 7886 11353 7903
rect 11336 7852 11353 7869
rect 11380 8022 11397 8039
rect 11380 7988 11397 8005
rect 11380 7954 11397 7971
rect 11380 7920 11397 7937
rect 11380 7886 11397 7903
rect 11380 7852 11397 7869
rect 11424 8022 11441 8039
rect 11424 7988 11441 8005
rect 11424 7954 11441 7971
rect 11424 7920 11441 7937
rect 11424 7886 11441 7903
rect 11424 7852 11441 7869
rect 11947 8022 11964 8039
rect 11947 7988 11964 8005
rect 11947 7954 11964 7971
rect 11947 7920 11964 7937
rect 11947 7886 11964 7903
rect 11947 7852 11964 7869
rect 11991 8022 12008 8039
rect 11991 7988 12008 8005
rect 11991 7954 12008 7971
rect 11991 7920 12008 7937
rect 11991 7886 12008 7903
rect 11991 7852 12008 7869
rect 12035 8022 12052 8039
rect 12035 7988 12052 8005
rect 12035 7954 12052 7971
rect 12035 7920 12052 7937
rect 12035 7886 12052 7903
rect 12035 7852 12052 7869
rect 12558 8022 12575 8039
rect 12558 7988 12575 8005
rect 12558 7954 12575 7971
rect 12558 7920 12575 7937
rect 12558 7886 12575 7903
rect 12558 7852 12575 7869
rect 12602 8022 12619 8039
rect 12602 7988 12619 8005
rect 12602 7954 12619 7971
rect 12602 7920 12619 7937
rect 12602 7886 12619 7903
rect 12602 7852 12619 7869
rect 12646 8022 12663 8039
rect 12646 7988 12663 8005
rect 12646 7954 12663 7971
rect 12646 7920 12663 7937
rect 12646 7886 12663 7903
rect 12646 7852 12663 7869
rect 9536 7372 9553 7389
rect 9536 7338 9553 7355
rect 9536 7304 9553 7321
rect 9536 7270 9553 7287
rect 9536 7236 9553 7253
rect 9536 7202 9553 7219
rect 9580 7372 9597 7389
rect 9580 7338 9597 7355
rect 9580 7304 9597 7321
rect 9580 7270 9597 7287
rect 9580 7236 9597 7253
rect 9580 7202 9597 7219
rect 9624 7372 9641 7389
rect 9624 7338 9641 7355
rect 9624 7304 9641 7321
rect 9624 7270 9641 7287
rect 9624 7236 9641 7253
rect 9624 7202 9641 7219
rect 10147 7372 10164 7389
rect 10147 7338 10164 7355
rect 10147 7304 10164 7321
rect 10147 7270 10164 7287
rect 10147 7236 10164 7253
rect 10147 7202 10164 7219
rect 10191 7372 10208 7389
rect 10191 7338 10208 7355
rect 10191 7304 10208 7321
rect 10191 7270 10208 7287
rect 10191 7236 10208 7253
rect 10191 7202 10208 7219
rect 10235 7372 10252 7389
rect 10235 7338 10252 7355
rect 10235 7304 10252 7321
rect 10235 7270 10252 7287
rect 10235 7236 10252 7253
rect 10235 7202 10252 7219
rect 10758 7372 10775 7389
rect 10758 7338 10775 7355
rect 10758 7304 10775 7321
rect 10758 7270 10775 7287
rect 10758 7236 10775 7253
rect 10758 7202 10775 7219
rect 10802 7372 10819 7389
rect 10802 7338 10819 7355
rect 10802 7304 10819 7321
rect 10802 7270 10819 7287
rect 10802 7236 10819 7253
rect 10802 7202 10819 7219
rect 10846 7372 10863 7389
rect 10846 7338 10863 7355
rect 10846 7304 10863 7321
rect 10846 7270 10863 7287
rect 10846 7236 10863 7253
rect 10846 7202 10863 7219
rect 11336 7372 11353 7389
rect 11336 7338 11353 7355
rect 11336 7304 11353 7321
rect 11336 7270 11353 7287
rect 11336 7236 11353 7253
rect 11336 7202 11353 7219
rect 11380 7372 11397 7389
rect 11380 7338 11397 7355
rect 11380 7304 11397 7321
rect 11380 7270 11397 7287
rect 11380 7236 11397 7253
rect 11380 7202 11397 7219
rect 11424 7372 11441 7389
rect 11424 7338 11441 7355
rect 11424 7304 11441 7321
rect 11424 7270 11441 7287
rect 11424 7236 11441 7253
rect 11424 7202 11441 7219
rect 11947 7372 11964 7389
rect 11947 7338 11964 7355
rect 11947 7304 11964 7321
rect 11947 7270 11964 7287
rect 11947 7236 11964 7253
rect 11947 7202 11964 7219
rect 11991 7372 12008 7389
rect 11991 7338 12008 7355
rect 11991 7304 12008 7321
rect 11991 7270 12008 7287
rect 11991 7236 12008 7253
rect 11991 7202 12008 7219
rect 12035 7372 12052 7389
rect 12035 7338 12052 7355
rect 12035 7304 12052 7321
rect 12035 7270 12052 7287
rect 12035 7236 12052 7253
rect 12035 7202 12052 7219
rect 12558 7372 12575 7389
rect 12558 7338 12575 7355
rect 12558 7304 12575 7321
rect 12558 7270 12575 7287
rect 12558 7236 12575 7253
rect 12558 7202 12575 7219
rect 12602 7372 12619 7389
rect 12602 7338 12619 7355
rect 12602 7304 12619 7321
rect 12602 7270 12619 7287
rect 12602 7236 12619 7253
rect 12602 7202 12619 7219
rect 12646 7372 12663 7389
rect 12646 7338 12663 7355
rect 12646 7304 12663 7321
rect 12646 7270 12663 7287
rect 12646 7236 12663 7253
rect 12646 7202 12663 7219
rect 9536 6732 9553 6749
rect 9536 6698 9553 6715
rect 9536 6664 9553 6681
rect 9536 6630 9553 6647
rect 9536 6596 9553 6613
rect 9536 6562 9553 6579
rect 9580 6732 9597 6749
rect 9580 6698 9597 6715
rect 9580 6664 9597 6681
rect 9580 6630 9597 6647
rect 9580 6596 9597 6613
rect 9580 6562 9597 6579
rect 9624 6732 9641 6749
rect 9624 6698 9641 6715
rect 9624 6664 9641 6681
rect 9624 6630 9641 6647
rect 9624 6596 9641 6613
rect 9624 6562 9641 6579
rect 10147 6732 10164 6749
rect 10147 6698 10164 6715
rect 10147 6664 10164 6681
rect 10147 6630 10164 6647
rect 10147 6596 10164 6613
rect 10147 6562 10164 6579
rect 10191 6732 10208 6749
rect 10191 6698 10208 6715
rect 10191 6664 10208 6681
rect 10191 6630 10208 6647
rect 10191 6596 10208 6613
rect 10191 6562 10208 6579
rect 10235 6732 10252 6749
rect 10235 6698 10252 6715
rect 10235 6664 10252 6681
rect 10235 6630 10252 6647
rect 10235 6596 10252 6613
rect 10235 6562 10252 6579
rect 10758 6732 10775 6749
rect 10758 6698 10775 6715
rect 10758 6664 10775 6681
rect 10758 6630 10775 6647
rect 10758 6596 10775 6613
rect 10758 6562 10775 6579
rect 10802 6732 10819 6749
rect 10802 6698 10819 6715
rect 10802 6664 10819 6681
rect 10802 6630 10819 6647
rect 10802 6596 10819 6613
rect 10802 6562 10819 6579
rect 10846 6732 10863 6749
rect 10846 6698 10863 6715
rect 10846 6664 10863 6681
rect 10846 6630 10863 6647
rect 10846 6596 10863 6613
rect 10846 6562 10863 6579
rect 11336 6732 11353 6749
rect 11336 6698 11353 6715
rect 11336 6664 11353 6681
rect 11336 6630 11353 6647
rect 11336 6596 11353 6613
rect 11336 6562 11353 6579
rect 11380 6732 11397 6749
rect 11380 6698 11397 6715
rect 11380 6664 11397 6681
rect 11380 6630 11397 6647
rect 11380 6596 11397 6613
rect 11380 6562 11397 6579
rect 11424 6732 11441 6749
rect 11424 6698 11441 6715
rect 11424 6664 11441 6681
rect 11424 6630 11441 6647
rect 11424 6596 11441 6613
rect 11424 6562 11441 6579
rect 11947 6732 11964 6749
rect 11947 6698 11964 6715
rect 11947 6664 11964 6681
rect 11947 6630 11964 6647
rect 11947 6596 11964 6613
rect 11947 6562 11964 6579
rect 11991 6732 12008 6749
rect 11991 6698 12008 6715
rect 11991 6664 12008 6681
rect 11991 6630 12008 6647
rect 11991 6596 12008 6613
rect 11991 6562 12008 6579
rect 12035 6732 12052 6749
rect 12035 6698 12052 6715
rect 12035 6664 12052 6681
rect 12035 6630 12052 6647
rect 12035 6596 12052 6613
rect 12035 6562 12052 6579
rect 12558 6732 12575 6749
rect 12558 6698 12575 6715
rect 12558 6664 12575 6681
rect 12558 6630 12575 6647
rect 12558 6596 12575 6613
rect 12558 6562 12575 6579
rect 12602 6732 12619 6749
rect 12602 6698 12619 6715
rect 12602 6664 12619 6681
rect 12602 6630 12619 6647
rect 12602 6596 12619 6613
rect 12602 6562 12619 6579
rect 12646 6732 12663 6749
rect 12646 6698 12663 6715
rect 12646 6664 12663 6681
rect 12646 6630 12663 6647
rect 12646 6596 12663 6613
rect 12646 6562 12663 6579
rect 9536 6082 9553 6099
rect 9536 6048 9553 6065
rect 9536 6014 9553 6031
rect 9536 5980 9553 5997
rect 9536 5946 9553 5963
rect 9536 5912 9553 5929
rect 9580 6082 9597 6099
rect 9580 6048 9597 6065
rect 9580 6014 9597 6031
rect 9580 5980 9597 5997
rect 9580 5946 9597 5963
rect 9580 5912 9597 5929
rect 9624 6082 9641 6099
rect 9624 6048 9641 6065
rect 9624 6014 9641 6031
rect 9624 5980 9641 5997
rect 9624 5946 9641 5963
rect 9624 5912 9641 5929
rect 10147 6082 10164 6099
rect 10147 6048 10164 6065
rect 10147 6014 10164 6031
rect 10147 5980 10164 5997
rect 10147 5946 10164 5963
rect 10147 5912 10164 5929
rect 10191 6082 10208 6099
rect 10191 6048 10208 6065
rect 10191 6014 10208 6031
rect 10191 5980 10208 5997
rect 10191 5946 10208 5963
rect 10191 5912 10208 5929
rect 10235 6082 10252 6099
rect 10235 6048 10252 6065
rect 10235 6014 10252 6031
rect 10235 5980 10252 5997
rect 10235 5946 10252 5963
rect 10235 5912 10252 5929
rect 10758 6082 10775 6099
rect 10758 6048 10775 6065
rect 10758 6014 10775 6031
rect 10758 5980 10775 5997
rect 10758 5946 10775 5963
rect 10758 5912 10775 5929
rect 10802 6082 10819 6099
rect 10802 6048 10819 6065
rect 10802 6014 10819 6031
rect 10802 5980 10819 5997
rect 10802 5946 10819 5963
rect 10802 5912 10819 5929
rect 10846 6082 10863 6099
rect 10846 6048 10863 6065
rect 10846 6014 10863 6031
rect 10846 5980 10863 5997
rect 10846 5946 10863 5963
rect 10846 5912 10863 5929
rect 11336 6082 11353 6099
rect 11336 6048 11353 6065
rect 11336 6014 11353 6031
rect 11336 5980 11353 5997
rect 11336 5946 11353 5963
rect 11336 5912 11353 5929
rect 11380 6082 11397 6099
rect 11380 6048 11397 6065
rect 11380 6014 11397 6031
rect 11380 5980 11397 5997
rect 11380 5946 11397 5963
rect 11380 5912 11397 5929
rect 11424 6082 11441 6099
rect 11424 6048 11441 6065
rect 11424 6014 11441 6031
rect 11424 5980 11441 5997
rect 11424 5946 11441 5963
rect 11424 5912 11441 5929
rect 11947 6082 11964 6099
rect 11947 6048 11964 6065
rect 11947 6014 11964 6031
rect 11947 5980 11964 5997
rect 11947 5946 11964 5963
rect 11947 5912 11964 5929
rect 11991 6082 12008 6099
rect 11991 6048 12008 6065
rect 11991 6014 12008 6031
rect 11991 5980 12008 5997
rect 11991 5946 12008 5963
rect 11991 5912 12008 5929
rect 12035 6082 12052 6099
rect 12035 6048 12052 6065
rect 12035 6014 12052 6031
rect 12035 5980 12052 5997
rect 12035 5946 12052 5963
rect 12035 5912 12052 5929
rect 12558 6082 12575 6099
rect 12558 6048 12575 6065
rect 12558 6014 12575 6031
rect 12558 5980 12575 5997
rect 12558 5946 12575 5963
rect 12558 5912 12575 5929
rect 12602 6082 12619 6099
rect 12602 6048 12619 6065
rect 12602 6014 12619 6031
rect 12602 5980 12619 5997
rect 12602 5946 12619 5963
rect 12602 5912 12619 5929
rect 12646 6082 12663 6099
rect 12646 6048 12663 6065
rect 12646 6014 12663 6031
rect 12646 5980 12663 5997
rect 12646 5946 12663 5963
rect 12646 5912 12663 5929
rect 9536 5432 9553 5449
rect 9536 5398 9553 5415
rect 9536 5364 9553 5381
rect 9536 5330 9553 5347
rect 9536 5296 9553 5313
rect 9536 5262 9553 5279
rect 9580 5432 9597 5449
rect 9580 5398 9597 5415
rect 9580 5364 9597 5381
rect 9580 5330 9597 5347
rect 9580 5296 9597 5313
rect 9580 5262 9597 5279
rect 9624 5432 9641 5449
rect 9624 5398 9641 5415
rect 9624 5364 9641 5381
rect 9624 5330 9641 5347
rect 9624 5296 9641 5313
rect 9624 5262 9641 5279
rect 10147 5432 10164 5449
rect 10147 5398 10164 5415
rect 10147 5364 10164 5381
rect 10147 5330 10164 5347
rect 10147 5296 10164 5313
rect 10147 5262 10164 5279
rect 10191 5432 10208 5449
rect 10191 5398 10208 5415
rect 10191 5364 10208 5381
rect 10191 5330 10208 5347
rect 10191 5296 10208 5313
rect 10191 5262 10208 5279
rect 10235 5432 10252 5449
rect 10235 5398 10252 5415
rect 10235 5364 10252 5381
rect 10235 5330 10252 5347
rect 10235 5296 10252 5313
rect 10235 5262 10252 5279
rect 10758 5432 10775 5449
rect 10758 5398 10775 5415
rect 10758 5364 10775 5381
rect 10758 5330 10775 5347
rect 10758 5296 10775 5313
rect 10758 5262 10775 5279
rect 10802 5432 10819 5449
rect 10802 5398 10819 5415
rect 10802 5364 10819 5381
rect 10802 5330 10819 5347
rect 10802 5296 10819 5313
rect 10802 5262 10819 5279
rect 10846 5432 10863 5449
rect 10846 5398 10863 5415
rect 10846 5364 10863 5381
rect 10846 5330 10863 5347
rect 10846 5296 10863 5313
rect 10846 5262 10863 5279
rect 11336 5432 11353 5449
rect 11336 5398 11353 5415
rect 11336 5364 11353 5381
rect 11336 5330 11353 5347
rect 11336 5296 11353 5313
rect 11336 5262 11353 5279
rect 11380 5432 11397 5449
rect 11380 5398 11397 5415
rect 11380 5364 11397 5381
rect 11380 5330 11397 5347
rect 11380 5296 11397 5313
rect 11380 5262 11397 5279
rect 11424 5432 11441 5449
rect 11424 5398 11441 5415
rect 11424 5364 11441 5381
rect 11424 5330 11441 5347
rect 11424 5296 11441 5313
rect 11424 5262 11441 5279
rect 11947 5432 11964 5449
rect 11947 5398 11964 5415
rect 11947 5364 11964 5381
rect 11947 5330 11964 5347
rect 11947 5296 11964 5313
rect 11947 5262 11964 5279
rect 11991 5432 12008 5449
rect 11991 5398 12008 5415
rect 11991 5364 12008 5381
rect 11991 5330 12008 5347
rect 11991 5296 12008 5313
rect 11991 5262 12008 5279
rect 12035 5432 12052 5449
rect 12035 5398 12052 5415
rect 12035 5364 12052 5381
rect 12035 5330 12052 5347
rect 12035 5296 12052 5313
rect 12035 5262 12052 5279
rect 12558 5432 12575 5449
rect 12558 5398 12575 5415
rect 12558 5364 12575 5381
rect 12558 5330 12575 5347
rect 12558 5296 12575 5313
rect 12558 5262 12575 5279
rect 12602 5432 12619 5449
rect 12602 5398 12619 5415
rect 12602 5364 12619 5381
rect 12602 5330 12619 5347
rect 12602 5296 12619 5313
rect 12602 5262 12619 5279
rect 12646 5432 12663 5449
rect 12646 5398 12663 5415
rect 12646 5364 12663 5381
rect 12646 5330 12663 5347
rect 12646 5296 12663 5313
rect 12646 5262 12663 5279
rect 9536 4792 9553 4809
rect 9536 4758 9553 4775
rect 9536 4724 9553 4741
rect 9536 4690 9553 4707
rect 9536 4656 9553 4673
rect 9536 4622 9553 4639
rect 9580 4792 9597 4809
rect 9580 4758 9597 4775
rect 9580 4724 9597 4741
rect 9580 4690 9597 4707
rect 9580 4656 9597 4673
rect 9580 4622 9597 4639
rect 9624 4792 9641 4809
rect 9624 4758 9641 4775
rect 9624 4724 9641 4741
rect 9624 4690 9641 4707
rect 9624 4656 9641 4673
rect 9624 4622 9641 4639
rect 10147 4792 10164 4809
rect 10147 4758 10164 4775
rect 10147 4724 10164 4741
rect 10147 4690 10164 4707
rect 10147 4656 10164 4673
rect 10147 4622 10164 4639
rect 10191 4792 10208 4809
rect 10191 4758 10208 4775
rect 10191 4724 10208 4741
rect 10191 4690 10208 4707
rect 10191 4656 10208 4673
rect 10191 4622 10208 4639
rect 10235 4792 10252 4809
rect 10235 4758 10252 4775
rect 10235 4724 10252 4741
rect 10235 4690 10252 4707
rect 10235 4656 10252 4673
rect 10235 4622 10252 4639
rect 10758 4792 10775 4809
rect 10758 4758 10775 4775
rect 10758 4724 10775 4741
rect 10758 4690 10775 4707
rect 10758 4656 10775 4673
rect 10758 4622 10775 4639
rect 10802 4792 10819 4809
rect 10802 4758 10819 4775
rect 10802 4724 10819 4741
rect 10802 4690 10819 4707
rect 10802 4656 10819 4673
rect 10802 4622 10819 4639
rect 10846 4792 10863 4809
rect 10846 4758 10863 4775
rect 10846 4724 10863 4741
rect 10846 4690 10863 4707
rect 10846 4656 10863 4673
rect 10846 4622 10863 4639
rect 11336 4792 11353 4809
rect 11336 4758 11353 4775
rect 11336 4724 11353 4741
rect 11336 4690 11353 4707
rect 11336 4656 11353 4673
rect 11336 4622 11353 4639
rect 11380 4792 11397 4809
rect 11380 4758 11397 4775
rect 11380 4724 11397 4741
rect 11380 4690 11397 4707
rect 11380 4656 11397 4673
rect 11380 4622 11397 4639
rect 11424 4792 11441 4809
rect 11424 4758 11441 4775
rect 11424 4724 11441 4741
rect 11424 4690 11441 4707
rect 11424 4656 11441 4673
rect 11424 4622 11441 4639
rect 11947 4792 11964 4809
rect 11947 4758 11964 4775
rect 11947 4724 11964 4741
rect 11947 4690 11964 4707
rect 11947 4656 11964 4673
rect 11947 4622 11964 4639
rect 11991 4792 12008 4809
rect 11991 4758 12008 4775
rect 11991 4724 12008 4741
rect 11991 4690 12008 4707
rect 11991 4656 12008 4673
rect 11991 4622 12008 4639
rect 12035 4792 12052 4809
rect 12035 4758 12052 4775
rect 12035 4724 12052 4741
rect 12035 4690 12052 4707
rect 12035 4656 12052 4673
rect 12035 4622 12052 4639
rect 12558 4792 12575 4809
rect 12558 4758 12575 4775
rect 12558 4724 12575 4741
rect 12558 4690 12575 4707
rect 12558 4656 12575 4673
rect 12558 4622 12575 4639
rect 12602 4792 12619 4809
rect 12602 4758 12619 4775
rect 12602 4724 12619 4741
rect 12602 4690 12619 4707
rect 12602 4656 12619 4673
rect 12602 4622 12619 4639
rect 12646 4792 12663 4809
rect 12646 4758 12663 4775
rect 12646 4724 12663 4741
rect 12646 4690 12663 4707
rect 12646 4656 12663 4673
rect 12646 4622 12663 4639
<< poly >>
rect 10170 8044 10185 8057
rect 10214 8044 10229 8057
rect 10781 8044 10796 8057
rect 10825 8044 10840 8057
rect 11359 8044 11374 8057
rect 11403 8044 11418 8057
rect 11970 8044 11985 8057
rect 12014 8044 12029 8057
rect 12581 8044 12596 8057
rect 12625 8044 12640 8057
rect 10170 7827 10185 7844
rect 10160 7819 10193 7827
rect 10160 7802 10168 7819
rect 10185 7802 10193 7819
rect 10160 7794 10193 7802
rect 10061 7767 10094 7775
rect 10061 7750 10069 7767
rect 10086 7757 10094 7767
rect 10086 7750 10141 7757
rect 10061 7742 10141 7750
rect 10061 7713 10105 7721
rect 10061 7696 10069 7713
rect 10086 7696 10105 7713
rect 10061 7688 10105 7696
rect 10090 7670 10105 7688
rect 10126 7670 10141 7742
rect 10170 7670 10185 7794
rect 10214 7773 10229 7844
rect 10781 7827 10796 7844
rect 10771 7819 10804 7827
rect 10771 7802 10779 7819
rect 10796 7802 10804 7819
rect 10771 7794 10804 7802
rect 10206 7765 10239 7773
rect 10206 7748 10214 7765
rect 10231 7748 10239 7765
rect 10206 7740 10239 7748
rect 10672 7767 10705 7775
rect 10672 7750 10680 7767
rect 10697 7757 10705 7767
rect 10697 7750 10752 7757
rect 10672 7742 10752 7750
rect 10214 7670 10229 7740
rect 10305 7729 10338 7737
rect 10305 7719 10313 7729
rect 10258 7712 10313 7719
rect 10330 7712 10338 7729
rect 10258 7704 10338 7712
rect 10672 7713 10716 7721
rect 10258 7670 10273 7704
rect 10672 7696 10680 7713
rect 10697 7696 10716 7713
rect 10672 7688 10716 7696
rect 10294 7670 10309 7683
rect 10701 7670 10716 7688
rect 10737 7670 10752 7742
rect 10781 7670 10796 7794
rect 10825 7773 10840 7844
rect 11359 7827 11374 7844
rect 11349 7819 11382 7827
rect 11349 7802 11357 7819
rect 11374 7802 11382 7819
rect 11349 7794 11382 7802
rect 10817 7765 10850 7773
rect 10817 7748 10825 7765
rect 10842 7748 10850 7765
rect 10817 7740 10850 7748
rect 11250 7767 11283 7775
rect 11250 7750 11258 7767
rect 11275 7757 11283 7767
rect 11275 7750 11330 7757
rect 11250 7742 11330 7750
rect 10825 7670 10840 7740
rect 10916 7729 10949 7737
rect 10916 7719 10924 7729
rect 10869 7712 10924 7719
rect 10941 7712 10949 7729
rect 10869 7704 10949 7712
rect 11250 7713 11294 7721
rect 10869 7670 10884 7704
rect 11250 7696 11258 7713
rect 11275 7696 11294 7713
rect 11250 7688 11294 7696
rect 10905 7670 10920 7683
rect 11279 7670 11294 7688
rect 11315 7670 11330 7742
rect 11359 7670 11374 7794
rect 11403 7773 11418 7844
rect 11970 7827 11985 7844
rect 11960 7819 11993 7827
rect 11960 7802 11968 7819
rect 11985 7802 11993 7819
rect 11960 7794 11993 7802
rect 11395 7765 11428 7773
rect 11395 7748 11403 7765
rect 11420 7748 11428 7765
rect 11395 7740 11428 7748
rect 11861 7767 11894 7775
rect 11861 7750 11869 7767
rect 11886 7757 11894 7767
rect 11886 7750 11941 7757
rect 11861 7742 11941 7750
rect 11403 7670 11418 7740
rect 11494 7729 11527 7737
rect 11494 7719 11502 7729
rect 11447 7712 11502 7719
rect 11519 7712 11527 7729
rect 11447 7704 11527 7712
rect 11861 7713 11905 7721
rect 11447 7670 11462 7704
rect 11861 7696 11869 7713
rect 11886 7696 11905 7713
rect 11861 7688 11905 7696
rect 11483 7670 11498 7683
rect 11890 7670 11905 7688
rect 11926 7670 11941 7742
rect 11970 7670 11985 7794
rect 12014 7773 12029 7844
rect 12581 7827 12596 7844
rect 12571 7819 12604 7827
rect 12571 7802 12579 7819
rect 12596 7802 12604 7819
rect 12571 7794 12604 7802
rect 12006 7765 12039 7773
rect 12006 7748 12014 7765
rect 12031 7748 12039 7765
rect 12006 7740 12039 7748
rect 12472 7767 12505 7775
rect 12472 7750 12480 7767
rect 12497 7757 12505 7767
rect 12497 7750 12552 7757
rect 12472 7742 12552 7750
rect 12014 7670 12029 7740
rect 12105 7729 12138 7737
rect 12105 7719 12113 7729
rect 12058 7712 12113 7719
rect 12130 7712 12138 7729
rect 12058 7704 12138 7712
rect 12472 7713 12516 7721
rect 12058 7670 12073 7704
rect 12472 7696 12480 7713
rect 12497 7696 12516 7713
rect 12472 7688 12516 7696
rect 12094 7670 12109 7683
rect 12501 7670 12516 7688
rect 12537 7670 12552 7742
rect 12581 7670 12596 7794
rect 12625 7773 12640 7844
rect 12617 7765 12650 7773
rect 12617 7748 12625 7765
rect 12642 7748 12650 7765
rect 12617 7740 12650 7748
rect 12625 7670 12640 7740
rect 12716 7729 12749 7737
rect 12716 7719 12724 7729
rect 12669 7712 12724 7719
rect 12741 7712 12749 7729
rect 12669 7704 12749 7712
rect 12669 7670 12684 7704
rect 12705 7670 12720 7683
rect 10090 7536 10105 7570
rect 10126 7557 10141 7570
rect 10170 7557 10185 7570
rect 10214 7557 10229 7570
rect 10258 7557 10273 7570
rect 10294 7536 10309 7570
rect 10090 7521 10309 7536
rect 10701 7536 10716 7570
rect 10737 7557 10752 7570
rect 10781 7557 10796 7570
rect 10825 7557 10840 7570
rect 10869 7557 10884 7570
rect 10905 7536 10920 7570
rect 10701 7521 10920 7536
rect 11279 7536 11294 7570
rect 11315 7557 11330 7570
rect 11359 7557 11374 7570
rect 11403 7557 11418 7570
rect 11447 7557 11462 7570
rect 11483 7536 11498 7570
rect 11279 7521 11498 7536
rect 11890 7536 11905 7570
rect 11926 7557 11941 7570
rect 11970 7557 11985 7570
rect 12014 7557 12029 7570
rect 12058 7557 12073 7570
rect 12094 7536 12109 7570
rect 11890 7521 12109 7536
rect 12501 7536 12516 7570
rect 12537 7557 12552 7570
rect 12581 7557 12596 7570
rect 12625 7557 12640 7570
rect 12669 7557 12684 7570
rect 12705 7536 12720 7570
rect 12501 7521 12720 7536
rect 9559 7394 9574 7407
rect 9603 7394 9618 7407
rect 10170 7394 10185 7407
rect 10214 7394 10229 7407
rect 10781 7394 10796 7407
rect 10825 7394 10840 7407
rect 11359 7394 11374 7407
rect 11403 7394 11418 7407
rect 11970 7394 11985 7407
rect 12014 7394 12029 7407
rect 12581 7394 12596 7407
rect 12625 7394 12640 7407
rect 9559 7177 9574 7194
rect 9549 7169 9582 7177
rect 9549 7152 9557 7169
rect 9574 7152 9582 7169
rect 9549 7144 9582 7152
rect 9450 7117 9483 7125
rect 9450 7100 9458 7117
rect 9475 7107 9483 7117
rect 9475 7100 9530 7107
rect 9450 7092 9530 7100
rect 9450 7063 9494 7071
rect 9450 7046 9458 7063
rect 9475 7046 9494 7063
rect 9450 7038 9494 7046
rect 9479 7020 9494 7038
rect 9515 7020 9530 7092
rect 9559 7020 9574 7144
rect 9603 7123 9618 7194
rect 10170 7177 10185 7194
rect 10160 7169 10193 7177
rect 10160 7152 10168 7169
rect 10185 7152 10193 7169
rect 10160 7144 10193 7152
rect 9595 7115 9628 7123
rect 9595 7098 9603 7115
rect 9620 7098 9628 7115
rect 9595 7090 9628 7098
rect 10061 7117 10094 7125
rect 10061 7100 10069 7117
rect 10086 7107 10094 7117
rect 10086 7100 10141 7107
rect 10061 7092 10141 7100
rect 9603 7020 9618 7090
rect 9694 7079 9727 7087
rect 9694 7069 9702 7079
rect 9647 7062 9702 7069
rect 9719 7062 9727 7079
rect 9647 7054 9727 7062
rect 10061 7063 10105 7071
rect 9647 7020 9662 7054
rect 10061 7046 10069 7063
rect 10086 7046 10105 7063
rect 10061 7038 10105 7046
rect 9683 7020 9698 7033
rect 10090 7020 10105 7038
rect 10126 7020 10141 7092
rect 10170 7020 10185 7144
rect 10214 7123 10229 7194
rect 10781 7177 10796 7194
rect 10771 7169 10804 7177
rect 10771 7152 10779 7169
rect 10796 7152 10804 7169
rect 10771 7144 10804 7152
rect 10206 7115 10239 7123
rect 10206 7098 10214 7115
rect 10231 7098 10239 7115
rect 10206 7090 10239 7098
rect 10672 7117 10705 7125
rect 10672 7100 10680 7117
rect 10697 7107 10705 7117
rect 10697 7100 10752 7107
rect 10672 7092 10752 7100
rect 10214 7020 10229 7090
rect 10305 7079 10338 7087
rect 10305 7069 10313 7079
rect 10258 7062 10313 7069
rect 10330 7062 10338 7079
rect 10258 7054 10338 7062
rect 10672 7063 10716 7071
rect 10258 7020 10273 7054
rect 10672 7046 10680 7063
rect 10697 7046 10716 7063
rect 10672 7038 10716 7046
rect 10294 7020 10309 7033
rect 10701 7020 10716 7038
rect 10737 7020 10752 7092
rect 10781 7020 10796 7144
rect 10825 7123 10840 7194
rect 11359 7177 11374 7194
rect 11349 7169 11382 7177
rect 11349 7152 11357 7169
rect 11374 7152 11382 7169
rect 11349 7144 11382 7152
rect 10817 7115 10850 7123
rect 10817 7098 10825 7115
rect 10842 7098 10850 7115
rect 10817 7090 10850 7098
rect 11250 7117 11283 7125
rect 11250 7100 11258 7117
rect 11275 7107 11283 7117
rect 11275 7100 11330 7107
rect 11250 7092 11330 7100
rect 10825 7020 10840 7090
rect 10916 7079 10949 7087
rect 10916 7069 10924 7079
rect 10869 7062 10924 7069
rect 10941 7062 10949 7079
rect 10869 7054 10949 7062
rect 11250 7063 11294 7071
rect 10869 7020 10884 7054
rect 11250 7046 11258 7063
rect 11275 7046 11294 7063
rect 11250 7038 11294 7046
rect 10905 7020 10920 7033
rect 11279 7020 11294 7038
rect 11315 7020 11330 7092
rect 11359 7020 11374 7144
rect 11403 7123 11418 7194
rect 11970 7177 11985 7194
rect 11960 7169 11993 7177
rect 11960 7152 11968 7169
rect 11985 7152 11993 7169
rect 11960 7144 11993 7152
rect 11395 7115 11428 7123
rect 11395 7098 11403 7115
rect 11420 7098 11428 7115
rect 11395 7090 11428 7098
rect 11861 7117 11894 7125
rect 11861 7100 11869 7117
rect 11886 7107 11894 7117
rect 11886 7100 11941 7107
rect 11861 7092 11941 7100
rect 11403 7020 11418 7090
rect 11494 7079 11527 7087
rect 11494 7069 11502 7079
rect 11447 7062 11502 7069
rect 11519 7062 11527 7079
rect 11447 7054 11527 7062
rect 11861 7063 11905 7071
rect 11447 7020 11462 7054
rect 11861 7046 11869 7063
rect 11886 7046 11905 7063
rect 11861 7038 11905 7046
rect 11483 7020 11498 7033
rect 11890 7020 11905 7038
rect 11926 7020 11941 7092
rect 11970 7020 11985 7144
rect 12014 7123 12029 7194
rect 12581 7177 12596 7194
rect 12571 7169 12604 7177
rect 12571 7152 12579 7169
rect 12596 7152 12604 7169
rect 12571 7144 12604 7152
rect 12006 7115 12039 7123
rect 12006 7098 12014 7115
rect 12031 7098 12039 7115
rect 12006 7090 12039 7098
rect 12472 7117 12505 7125
rect 12472 7100 12480 7117
rect 12497 7107 12505 7117
rect 12497 7100 12552 7107
rect 12472 7092 12552 7100
rect 12014 7020 12029 7090
rect 12105 7079 12138 7087
rect 12105 7069 12113 7079
rect 12058 7062 12113 7069
rect 12130 7062 12138 7079
rect 12058 7054 12138 7062
rect 12472 7063 12516 7071
rect 12058 7020 12073 7054
rect 12472 7046 12480 7063
rect 12497 7046 12516 7063
rect 12472 7038 12516 7046
rect 12094 7020 12109 7033
rect 12501 7020 12516 7038
rect 12537 7020 12552 7092
rect 12581 7020 12596 7144
rect 12625 7123 12640 7194
rect 12617 7115 12650 7123
rect 12617 7098 12625 7115
rect 12642 7098 12650 7115
rect 12617 7090 12650 7098
rect 12625 7020 12640 7090
rect 12716 7079 12749 7087
rect 12716 7069 12724 7079
rect 12669 7062 12724 7069
rect 12741 7062 12749 7079
rect 12669 7054 12749 7062
rect 12669 7020 12684 7054
rect 12705 7020 12720 7033
rect 9479 6886 9494 6920
rect 9515 6907 9530 6920
rect 9559 6907 9574 6920
rect 9603 6907 9618 6920
rect 9647 6907 9662 6920
rect 9683 6886 9698 6920
rect 9479 6871 9698 6886
rect 10090 6886 10105 6920
rect 10126 6907 10141 6920
rect 10170 6907 10185 6920
rect 10214 6907 10229 6920
rect 10258 6907 10273 6920
rect 10294 6886 10309 6920
rect 10090 6871 10309 6886
rect 10701 6886 10716 6920
rect 10737 6907 10752 6920
rect 10781 6907 10796 6920
rect 10825 6907 10840 6920
rect 10869 6907 10884 6920
rect 10905 6886 10920 6920
rect 10701 6871 10920 6886
rect 11279 6886 11294 6920
rect 11315 6907 11330 6920
rect 11359 6907 11374 6920
rect 11403 6907 11418 6920
rect 11447 6907 11462 6920
rect 11483 6886 11498 6920
rect 11279 6871 11498 6886
rect 11890 6886 11905 6920
rect 11926 6907 11941 6920
rect 11970 6907 11985 6920
rect 12014 6907 12029 6920
rect 12058 6907 12073 6920
rect 12094 6886 12109 6920
rect 11890 6871 12109 6886
rect 12501 6886 12516 6920
rect 12537 6907 12552 6920
rect 12581 6907 12596 6920
rect 12625 6907 12640 6920
rect 12669 6907 12684 6920
rect 12705 6886 12720 6920
rect 12501 6871 12720 6886
rect 9559 6754 9574 6767
rect 9603 6754 9618 6767
rect 10170 6754 10185 6767
rect 10214 6754 10229 6767
rect 10781 6754 10796 6767
rect 10825 6754 10840 6767
rect 11359 6754 11374 6767
rect 11403 6754 11418 6767
rect 11970 6754 11985 6767
rect 12014 6754 12029 6767
rect 12581 6754 12596 6767
rect 12625 6754 12640 6767
rect 9559 6537 9574 6554
rect 9549 6529 9582 6537
rect 9549 6512 9557 6529
rect 9574 6512 9582 6529
rect 9549 6504 9582 6512
rect 9450 6477 9483 6485
rect 9450 6460 9458 6477
rect 9475 6467 9483 6477
rect 9475 6460 9530 6467
rect 9450 6452 9530 6460
rect 9450 6423 9494 6431
rect 9450 6406 9458 6423
rect 9475 6406 9494 6423
rect 9450 6398 9494 6406
rect 9479 6380 9494 6398
rect 9515 6380 9530 6452
rect 9559 6380 9574 6504
rect 9603 6483 9618 6554
rect 10170 6537 10185 6554
rect 10160 6529 10193 6537
rect 10160 6512 10168 6529
rect 10185 6512 10193 6529
rect 10160 6504 10193 6512
rect 9595 6475 9628 6483
rect 9595 6458 9603 6475
rect 9620 6458 9628 6475
rect 9595 6450 9628 6458
rect 10061 6477 10094 6485
rect 10061 6460 10069 6477
rect 10086 6467 10094 6477
rect 10086 6460 10141 6467
rect 10061 6452 10141 6460
rect 9603 6380 9618 6450
rect 9694 6439 9727 6447
rect 9694 6429 9702 6439
rect 9647 6422 9702 6429
rect 9719 6422 9727 6439
rect 9647 6414 9727 6422
rect 10061 6423 10105 6431
rect 9647 6380 9662 6414
rect 10061 6406 10069 6423
rect 10086 6406 10105 6423
rect 10061 6398 10105 6406
rect 9683 6380 9698 6393
rect 10090 6380 10105 6398
rect 10126 6380 10141 6452
rect 10170 6380 10185 6504
rect 10214 6483 10229 6554
rect 10781 6537 10796 6554
rect 10771 6529 10804 6537
rect 10771 6512 10779 6529
rect 10796 6512 10804 6529
rect 10771 6504 10804 6512
rect 10206 6475 10239 6483
rect 10206 6458 10214 6475
rect 10231 6458 10239 6475
rect 10206 6450 10239 6458
rect 10672 6477 10705 6485
rect 10672 6460 10680 6477
rect 10697 6467 10705 6477
rect 10697 6460 10752 6467
rect 10672 6452 10752 6460
rect 10214 6380 10229 6450
rect 10305 6439 10338 6447
rect 10305 6429 10313 6439
rect 10258 6422 10313 6429
rect 10330 6422 10338 6439
rect 10258 6414 10338 6422
rect 10672 6423 10716 6431
rect 10258 6380 10273 6414
rect 10672 6406 10680 6423
rect 10697 6406 10716 6423
rect 10672 6398 10716 6406
rect 10294 6380 10309 6393
rect 10701 6380 10716 6398
rect 10737 6380 10752 6452
rect 10781 6380 10796 6504
rect 10825 6483 10840 6554
rect 11359 6537 11374 6554
rect 11349 6529 11382 6537
rect 11349 6512 11357 6529
rect 11374 6512 11382 6529
rect 11349 6504 11382 6512
rect 10817 6475 10850 6483
rect 10817 6458 10825 6475
rect 10842 6458 10850 6475
rect 10817 6450 10850 6458
rect 11250 6477 11283 6485
rect 11250 6460 11258 6477
rect 11275 6467 11283 6477
rect 11275 6460 11330 6467
rect 11250 6452 11330 6460
rect 10825 6380 10840 6450
rect 10916 6439 10949 6447
rect 10916 6429 10924 6439
rect 10869 6422 10924 6429
rect 10941 6422 10949 6439
rect 10869 6414 10949 6422
rect 11250 6423 11294 6431
rect 10869 6380 10884 6414
rect 11250 6406 11258 6423
rect 11275 6406 11294 6423
rect 11250 6398 11294 6406
rect 10905 6380 10920 6393
rect 11279 6380 11294 6398
rect 11315 6380 11330 6452
rect 11359 6380 11374 6504
rect 11403 6483 11418 6554
rect 11970 6537 11985 6554
rect 11960 6529 11993 6537
rect 11960 6512 11968 6529
rect 11985 6512 11993 6529
rect 11960 6504 11993 6512
rect 11395 6475 11428 6483
rect 11395 6458 11403 6475
rect 11420 6458 11428 6475
rect 11395 6450 11428 6458
rect 11861 6477 11894 6485
rect 11861 6460 11869 6477
rect 11886 6467 11894 6477
rect 11886 6460 11941 6467
rect 11861 6452 11941 6460
rect 11403 6380 11418 6450
rect 11494 6439 11527 6447
rect 11494 6429 11502 6439
rect 11447 6422 11502 6429
rect 11519 6422 11527 6439
rect 11447 6414 11527 6422
rect 11861 6423 11905 6431
rect 11447 6380 11462 6414
rect 11861 6406 11869 6423
rect 11886 6406 11905 6423
rect 11861 6398 11905 6406
rect 11483 6380 11498 6393
rect 11890 6380 11905 6398
rect 11926 6380 11941 6452
rect 11970 6380 11985 6504
rect 12014 6483 12029 6554
rect 12581 6537 12596 6554
rect 12571 6529 12604 6537
rect 12571 6512 12579 6529
rect 12596 6512 12604 6529
rect 12571 6504 12604 6512
rect 12006 6475 12039 6483
rect 12006 6458 12014 6475
rect 12031 6458 12039 6475
rect 12006 6450 12039 6458
rect 12472 6477 12505 6485
rect 12472 6460 12480 6477
rect 12497 6467 12505 6477
rect 12497 6460 12552 6467
rect 12472 6452 12552 6460
rect 12014 6380 12029 6450
rect 12105 6439 12138 6447
rect 12105 6429 12113 6439
rect 12058 6422 12113 6429
rect 12130 6422 12138 6439
rect 12058 6414 12138 6422
rect 12472 6423 12516 6431
rect 12058 6380 12073 6414
rect 12472 6406 12480 6423
rect 12497 6406 12516 6423
rect 12472 6398 12516 6406
rect 12094 6380 12109 6393
rect 12501 6380 12516 6398
rect 12537 6380 12552 6452
rect 12581 6380 12596 6504
rect 12625 6483 12640 6554
rect 12617 6475 12650 6483
rect 12617 6458 12625 6475
rect 12642 6458 12650 6475
rect 12617 6450 12650 6458
rect 12625 6380 12640 6450
rect 12716 6439 12749 6447
rect 12716 6429 12724 6439
rect 12669 6422 12724 6429
rect 12741 6422 12749 6439
rect 12669 6414 12749 6422
rect 12669 6380 12684 6414
rect 12705 6380 12720 6393
rect 9479 6246 9494 6280
rect 9515 6267 9530 6280
rect 9559 6267 9574 6280
rect 9603 6267 9618 6280
rect 9647 6267 9662 6280
rect 9683 6246 9698 6280
rect 9479 6231 9698 6246
rect 10090 6246 10105 6280
rect 10126 6267 10141 6280
rect 10170 6267 10185 6280
rect 10214 6267 10229 6280
rect 10258 6267 10273 6280
rect 10294 6246 10309 6280
rect 10090 6231 10309 6246
rect 10701 6246 10716 6280
rect 10737 6267 10752 6280
rect 10781 6267 10796 6280
rect 10825 6267 10840 6280
rect 10869 6267 10884 6280
rect 10905 6246 10920 6280
rect 10701 6231 10920 6246
rect 11279 6246 11294 6280
rect 11315 6267 11330 6280
rect 11359 6267 11374 6280
rect 11403 6267 11418 6280
rect 11447 6267 11462 6280
rect 11483 6246 11498 6280
rect 11279 6231 11498 6246
rect 11890 6246 11905 6280
rect 11926 6267 11941 6280
rect 11970 6267 11985 6280
rect 12014 6267 12029 6280
rect 12058 6267 12073 6280
rect 12094 6246 12109 6280
rect 11890 6231 12109 6246
rect 12501 6246 12516 6280
rect 12537 6267 12552 6280
rect 12581 6267 12596 6280
rect 12625 6267 12640 6280
rect 12669 6267 12684 6280
rect 12705 6246 12720 6280
rect 12501 6231 12720 6246
rect 9559 6104 9574 6117
rect 9603 6104 9618 6117
rect 10170 6104 10185 6117
rect 10214 6104 10229 6117
rect 10781 6104 10796 6117
rect 10825 6104 10840 6117
rect 11359 6104 11374 6117
rect 11403 6104 11418 6117
rect 11970 6104 11985 6117
rect 12014 6104 12029 6117
rect 12581 6104 12596 6117
rect 12625 6104 12640 6117
rect 9559 5887 9574 5904
rect 9549 5879 9582 5887
rect 9549 5862 9557 5879
rect 9574 5862 9582 5879
rect 9549 5854 9582 5862
rect 9450 5827 9483 5835
rect 9450 5810 9458 5827
rect 9475 5817 9483 5827
rect 9475 5810 9530 5817
rect 9450 5802 9530 5810
rect 9450 5773 9494 5781
rect 9450 5756 9458 5773
rect 9475 5756 9494 5773
rect 9450 5748 9494 5756
rect 9479 5730 9494 5748
rect 9515 5730 9530 5802
rect 9559 5730 9574 5854
rect 9603 5833 9618 5904
rect 10170 5887 10185 5904
rect 10160 5879 10193 5887
rect 10160 5862 10168 5879
rect 10185 5862 10193 5879
rect 10160 5854 10193 5862
rect 9595 5825 9628 5833
rect 9595 5808 9603 5825
rect 9620 5808 9628 5825
rect 9595 5800 9628 5808
rect 10061 5827 10094 5835
rect 10061 5810 10069 5827
rect 10086 5817 10094 5827
rect 10086 5810 10141 5817
rect 10061 5802 10141 5810
rect 9603 5730 9618 5800
rect 9694 5789 9727 5797
rect 9694 5779 9702 5789
rect 9647 5772 9702 5779
rect 9719 5772 9727 5789
rect 9647 5764 9727 5772
rect 10061 5773 10105 5781
rect 9647 5730 9662 5764
rect 10061 5756 10069 5773
rect 10086 5756 10105 5773
rect 10061 5748 10105 5756
rect 9683 5730 9698 5743
rect 10090 5730 10105 5748
rect 10126 5730 10141 5802
rect 10170 5730 10185 5854
rect 10214 5833 10229 5904
rect 10781 5887 10796 5904
rect 10771 5879 10804 5887
rect 10771 5862 10779 5879
rect 10796 5862 10804 5879
rect 10771 5854 10804 5862
rect 10206 5825 10239 5833
rect 10206 5808 10214 5825
rect 10231 5808 10239 5825
rect 10206 5800 10239 5808
rect 10672 5827 10705 5835
rect 10672 5810 10680 5827
rect 10697 5817 10705 5827
rect 10697 5810 10752 5817
rect 10672 5802 10752 5810
rect 10214 5730 10229 5800
rect 10305 5789 10338 5797
rect 10305 5779 10313 5789
rect 10258 5772 10313 5779
rect 10330 5772 10338 5789
rect 10258 5764 10338 5772
rect 10672 5773 10716 5781
rect 10258 5730 10273 5764
rect 10672 5756 10680 5773
rect 10697 5756 10716 5773
rect 10672 5748 10716 5756
rect 10294 5730 10309 5743
rect 10701 5730 10716 5748
rect 10737 5730 10752 5802
rect 10781 5730 10796 5854
rect 10825 5833 10840 5904
rect 11359 5887 11374 5904
rect 11349 5879 11382 5887
rect 11349 5862 11357 5879
rect 11374 5862 11382 5879
rect 11349 5854 11382 5862
rect 10817 5825 10850 5833
rect 10817 5808 10825 5825
rect 10842 5808 10850 5825
rect 10817 5800 10850 5808
rect 11250 5827 11283 5835
rect 11250 5810 11258 5827
rect 11275 5817 11283 5827
rect 11275 5810 11330 5817
rect 11250 5802 11330 5810
rect 10825 5730 10840 5800
rect 10916 5789 10949 5797
rect 10916 5779 10924 5789
rect 10869 5772 10924 5779
rect 10941 5772 10949 5789
rect 10869 5764 10949 5772
rect 11250 5773 11294 5781
rect 10869 5730 10884 5764
rect 11250 5756 11258 5773
rect 11275 5756 11294 5773
rect 11250 5748 11294 5756
rect 10905 5730 10920 5743
rect 11279 5730 11294 5748
rect 11315 5730 11330 5802
rect 11359 5730 11374 5854
rect 11403 5833 11418 5904
rect 11970 5887 11985 5904
rect 11960 5879 11993 5887
rect 11960 5862 11968 5879
rect 11985 5862 11993 5879
rect 11960 5854 11993 5862
rect 11395 5825 11428 5833
rect 11395 5808 11403 5825
rect 11420 5808 11428 5825
rect 11395 5800 11428 5808
rect 11861 5827 11894 5835
rect 11861 5810 11869 5827
rect 11886 5817 11894 5827
rect 11886 5810 11941 5817
rect 11861 5802 11941 5810
rect 11403 5730 11418 5800
rect 11494 5789 11527 5797
rect 11494 5779 11502 5789
rect 11447 5772 11502 5779
rect 11519 5772 11527 5789
rect 11447 5764 11527 5772
rect 11861 5773 11905 5781
rect 11447 5730 11462 5764
rect 11861 5756 11869 5773
rect 11886 5756 11905 5773
rect 11861 5748 11905 5756
rect 11483 5730 11498 5743
rect 11890 5730 11905 5748
rect 11926 5730 11941 5802
rect 11970 5730 11985 5854
rect 12014 5833 12029 5904
rect 12581 5887 12596 5904
rect 12571 5879 12604 5887
rect 12571 5862 12579 5879
rect 12596 5862 12604 5879
rect 12571 5854 12604 5862
rect 12006 5825 12039 5833
rect 12006 5808 12014 5825
rect 12031 5808 12039 5825
rect 12006 5800 12039 5808
rect 12472 5827 12505 5835
rect 12472 5810 12480 5827
rect 12497 5817 12505 5827
rect 12497 5810 12552 5817
rect 12472 5802 12552 5810
rect 12014 5730 12029 5800
rect 12105 5789 12138 5797
rect 12105 5779 12113 5789
rect 12058 5772 12113 5779
rect 12130 5772 12138 5789
rect 12058 5764 12138 5772
rect 12472 5773 12516 5781
rect 12058 5730 12073 5764
rect 12472 5756 12480 5773
rect 12497 5756 12516 5773
rect 12472 5748 12516 5756
rect 12094 5730 12109 5743
rect 12501 5730 12516 5748
rect 12537 5730 12552 5802
rect 12581 5730 12596 5854
rect 12625 5833 12640 5904
rect 12617 5825 12650 5833
rect 12617 5808 12625 5825
rect 12642 5808 12650 5825
rect 12617 5800 12650 5808
rect 12625 5730 12640 5800
rect 12716 5789 12749 5797
rect 12716 5779 12724 5789
rect 12669 5772 12724 5779
rect 12741 5772 12749 5789
rect 12669 5764 12749 5772
rect 12669 5730 12684 5764
rect 12705 5730 12720 5743
rect 9479 5596 9494 5630
rect 9515 5617 9530 5630
rect 9559 5617 9574 5630
rect 9603 5617 9618 5630
rect 9647 5617 9662 5630
rect 9683 5596 9698 5630
rect 9479 5581 9698 5596
rect 10090 5596 10105 5630
rect 10126 5617 10141 5630
rect 10170 5617 10185 5630
rect 10214 5617 10229 5630
rect 10258 5617 10273 5630
rect 10294 5596 10309 5630
rect 10090 5581 10309 5596
rect 10701 5596 10716 5630
rect 10737 5617 10752 5630
rect 10781 5617 10796 5630
rect 10825 5617 10840 5630
rect 10869 5617 10884 5630
rect 10905 5596 10920 5630
rect 10701 5581 10920 5596
rect 11279 5596 11294 5630
rect 11315 5617 11330 5630
rect 11359 5617 11374 5630
rect 11403 5617 11418 5630
rect 11447 5617 11462 5630
rect 11483 5596 11498 5630
rect 11279 5581 11498 5596
rect 11890 5596 11905 5630
rect 11926 5617 11941 5630
rect 11970 5617 11985 5630
rect 12014 5617 12029 5630
rect 12058 5617 12073 5630
rect 12094 5596 12109 5630
rect 11890 5581 12109 5596
rect 12501 5596 12516 5630
rect 12537 5617 12552 5630
rect 12581 5617 12596 5630
rect 12625 5617 12640 5630
rect 12669 5617 12684 5630
rect 12705 5596 12720 5630
rect 12501 5581 12720 5596
rect 9559 5454 9574 5467
rect 9603 5454 9618 5467
rect 10170 5454 10185 5467
rect 10214 5454 10229 5467
rect 10781 5454 10796 5467
rect 10825 5454 10840 5467
rect 11359 5454 11374 5467
rect 11403 5454 11418 5467
rect 11970 5454 11985 5467
rect 12014 5454 12029 5467
rect 12581 5454 12596 5467
rect 12625 5454 12640 5467
rect 9559 5237 9574 5254
rect 9549 5229 9582 5237
rect 9549 5212 9557 5229
rect 9574 5212 9582 5229
rect 9549 5204 9582 5212
rect 9450 5177 9483 5185
rect 9450 5160 9458 5177
rect 9475 5167 9483 5177
rect 9475 5160 9530 5167
rect 9450 5152 9530 5160
rect 9450 5123 9494 5131
rect 9450 5106 9458 5123
rect 9475 5106 9494 5123
rect 9450 5098 9494 5106
rect 9479 5080 9494 5098
rect 9515 5080 9530 5152
rect 9559 5080 9574 5204
rect 9603 5183 9618 5254
rect 10170 5237 10185 5254
rect 10160 5229 10193 5237
rect 10160 5212 10168 5229
rect 10185 5212 10193 5229
rect 10160 5204 10193 5212
rect 9595 5175 9628 5183
rect 9595 5158 9603 5175
rect 9620 5158 9628 5175
rect 9595 5150 9628 5158
rect 10061 5177 10094 5185
rect 10061 5160 10069 5177
rect 10086 5167 10094 5177
rect 10086 5160 10141 5167
rect 10061 5152 10141 5160
rect 9603 5080 9618 5150
rect 9694 5139 9727 5147
rect 9694 5129 9702 5139
rect 9647 5122 9702 5129
rect 9719 5122 9727 5139
rect 9647 5114 9727 5122
rect 10061 5123 10105 5131
rect 9647 5080 9662 5114
rect 10061 5106 10069 5123
rect 10086 5106 10105 5123
rect 10061 5098 10105 5106
rect 9683 5080 9698 5093
rect 10090 5080 10105 5098
rect 10126 5080 10141 5152
rect 10170 5080 10185 5204
rect 10214 5183 10229 5254
rect 10781 5237 10796 5254
rect 10771 5229 10804 5237
rect 10771 5212 10779 5229
rect 10796 5212 10804 5229
rect 10771 5204 10804 5212
rect 10206 5175 10239 5183
rect 10206 5158 10214 5175
rect 10231 5158 10239 5175
rect 10206 5150 10239 5158
rect 10672 5177 10705 5185
rect 10672 5160 10680 5177
rect 10697 5167 10705 5177
rect 10697 5160 10752 5167
rect 10672 5152 10752 5160
rect 10214 5080 10229 5150
rect 10305 5139 10338 5147
rect 10305 5129 10313 5139
rect 10258 5122 10313 5129
rect 10330 5122 10338 5139
rect 10258 5114 10338 5122
rect 10672 5123 10716 5131
rect 10258 5080 10273 5114
rect 10672 5106 10680 5123
rect 10697 5106 10716 5123
rect 10672 5098 10716 5106
rect 10294 5080 10309 5093
rect 10701 5080 10716 5098
rect 10737 5080 10752 5152
rect 10781 5080 10796 5204
rect 10825 5183 10840 5254
rect 11359 5237 11374 5254
rect 11349 5229 11382 5237
rect 11349 5212 11357 5229
rect 11374 5212 11382 5229
rect 11349 5204 11382 5212
rect 10817 5175 10850 5183
rect 10817 5158 10825 5175
rect 10842 5158 10850 5175
rect 10817 5150 10850 5158
rect 11250 5177 11283 5185
rect 11250 5160 11258 5177
rect 11275 5167 11283 5177
rect 11275 5160 11330 5167
rect 11250 5152 11330 5160
rect 10825 5080 10840 5150
rect 10916 5139 10949 5147
rect 10916 5129 10924 5139
rect 10869 5122 10924 5129
rect 10941 5122 10949 5139
rect 10869 5114 10949 5122
rect 11250 5123 11294 5131
rect 10869 5080 10884 5114
rect 11250 5106 11258 5123
rect 11275 5106 11294 5123
rect 11250 5098 11294 5106
rect 10905 5080 10920 5093
rect 11279 5080 11294 5098
rect 11315 5080 11330 5152
rect 11359 5080 11374 5204
rect 11403 5183 11418 5254
rect 11970 5237 11985 5254
rect 11960 5229 11993 5237
rect 11960 5212 11968 5229
rect 11985 5212 11993 5229
rect 11960 5204 11993 5212
rect 11395 5175 11428 5183
rect 11395 5158 11403 5175
rect 11420 5158 11428 5175
rect 11395 5150 11428 5158
rect 11861 5177 11894 5185
rect 11861 5160 11869 5177
rect 11886 5167 11894 5177
rect 11886 5160 11941 5167
rect 11861 5152 11941 5160
rect 11403 5080 11418 5150
rect 11494 5139 11527 5147
rect 11494 5129 11502 5139
rect 11447 5122 11502 5129
rect 11519 5122 11527 5139
rect 11447 5114 11527 5122
rect 11861 5123 11905 5131
rect 11447 5080 11462 5114
rect 11861 5106 11869 5123
rect 11886 5106 11905 5123
rect 11861 5098 11905 5106
rect 11483 5080 11498 5093
rect 11890 5080 11905 5098
rect 11926 5080 11941 5152
rect 11970 5080 11985 5204
rect 12014 5183 12029 5254
rect 12581 5237 12596 5254
rect 12571 5229 12604 5237
rect 12571 5212 12579 5229
rect 12596 5212 12604 5229
rect 12571 5204 12604 5212
rect 12006 5175 12039 5183
rect 12006 5158 12014 5175
rect 12031 5158 12039 5175
rect 12006 5150 12039 5158
rect 12472 5177 12505 5185
rect 12472 5160 12480 5177
rect 12497 5167 12505 5177
rect 12497 5160 12552 5167
rect 12472 5152 12552 5160
rect 12014 5080 12029 5150
rect 12105 5139 12138 5147
rect 12105 5129 12113 5139
rect 12058 5122 12113 5129
rect 12130 5122 12138 5139
rect 12058 5114 12138 5122
rect 12472 5123 12516 5131
rect 12058 5080 12073 5114
rect 12472 5106 12480 5123
rect 12497 5106 12516 5123
rect 12472 5098 12516 5106
rect 12094 5080 12109 5093
rect 12501 5080 12516 5098
rect 12537 5080 12552 5152
rect 12581 5080 12596 5204
rect 12625 5183 12640 5254
rect 12617 5175 12650 5183
rect 12617 5158 12625 5175
rect 12642 5158 12650 5175
rect 12617 5150 12650 5158
rect 12625 5080 12640 5150
rect 12716 5139 12749 5147
rect 12716 5129 12724 5139
rect 12669 5122 12724 5129
rect 12741 5122 12749 5139
rect 12669 5114 12749 5122
rect 12669 5080 12684 5114
rect 12705 5080 12720 5093
rect 9479 4946 9494 4980
rect 9515 4967 9530 4980
rect 9559 4967 9574 4980
rect 9603 4967 9618 4980
rect 9647 4967 9662 4980
rect 9683 4946 9698 4980
rect 9479 4931 9698 4946
rect 10090 4946 10105 4980
rect 10126 4967 10141 4980
rect 10170 4967 10185 4980
rect 10214 4967 10229 4980
rect 10258 4967 10273 4980
rect 10294 4946 10309 4980
rect 10090 4931 10309 4946
rect 10701 4946 10716 4980
rect 10737 4967 10752 4980
rect 10781 4967 10796 4980
rect 10825 4967 10840 4980
rect 10869 4967 10884 4980
rect 10905 4946 10920 4980
rect 10701 4931 10920 4946
rect 11279 4946 11294 4980
rect 11315 4967 11330 4980
rect 11359 4967 11374 4980
rect 11403 4967 11418 4980
rect 11447 4967 11462 4980
rect 11483 4946 11498 4980
rect 11279 4931 11498 4946
rect 11890 4946 11905 4980
rect 11926 4967 11941 4980
rect 11970 4967 11985 4980
rect 12014 4967 12029 4980
rect 12058 4967 12073 4980
rect 12094 4946 12109 4980
rect 11890 4931 12109 4946
rect 12501 4946 12516 4980
rect 12537 4967 12552 4980
rect 12581 4967 12596 4980
rect 12625 4967 12640 4980
rect 12669 4967 12684 4980
rect 12705 4946 12720 4980
rect 12501 4931 12720 4946
rect 9559 4814 9574 4827
rect 9603 4814 9618 4827
rect 10170 4814 10185 4827
rect 10214 4814 10229 4827
rect 10781 4814 10796 4827
rect 10825 4814 10840 4827
rect 11359 4814 11374 4827
rect 11403 4814 11418 4827
rect 11970 4814 11985 4827
rect 12014 4814 12029 4827
rect 12581 4814 12596 4827
rect 12625 4814 12640 4827
rect 9559 4597 9574 4614
rect 9549 4589 9582 4597
rect 9549 4572 9557 4589
rect 9574 4572 9582 4589
rect 9549 4564 9582 4572
rect 9450 4537 9483 4545
rect 9450 4520 9458 4537
rect 9475 4527 9483 4537
rect 9475 4520 9530 4527
rect 9450 4512 9530 4520
rect 9450 4483 9494 4491
rect 9450 4466 9458 4483
rect 9475 4466 9494 4483
rect 9450 4458 9494 4466
rect 9479 4440 9494 4458
rect 9515 4440 9530 4512
rect 9559 4440 9574 4564
rect 9603 4543 9618 4614
rect 10170 4597 10185 4614
rect 10160 4589 10193 4597
rect 10160 4572 10168 4589
rect 10185 4572 10193 4589
rect 10160 4564 10193 4572
rect 9595 4535 9628 4543
rect 9595 4518 9603 4535
rect 9620 4518 9628 4535
rect 9595 4510 9628 4518
rect 10061 4537 10094 4545
rect 10061 4520 10069 4537
rect 10086 4527 10094 4537
rect 10086 4520 10141 4527
rect 10061 4512 10141 4520
rect 9603 4440 9618 4510
rect 9694 4499 9727 4507
rect 9694 4489 9702 4499
rect 9647 4482 9702 4489
rect 9719 4482 9727 4499
rect 9647 4474 9727 4482
rect 10061 4483 10105 4491
rect 9647 4440 9662 4474
rect 10061 4466 10069 4483
rect 10086 4466 10105 4483
rect 10061 4458 10105 4466
rect 9683 4440 9698 4453
rect 10090 4440 10105 4458
rect 10126 4440 10141 4512
rect 10170 4440 10185 4564
rect 10214 4543 10229 4614
rect 10781 4597 10796 4614
rect 10771 4589 10804 4597
rect 10771 4572 10779 4589
rect 10796 4572 10804 4589
rect 10771 4564 10804 4572
rect 10206 4535 10239 4543
rect 10206 4518 10214 4535
rect 10231 4518 10239 4535
rect 10206 4510 10239 4518
rect 10672 4537 10705 4545
rect 10672 4520 10680 4537
rect 10697 4527 10705 4537
rect 10697 4520 10752 4527
rect 10672 4512 10752 4520
rect 10214 4440 10229 4510
rect 10305 4499 10338 4507
rect 10305 4489 10313 4499
rect 10258 4482 10313 4489
rect 10330 4482 10338 4499
rect 10258 4474 10338 4482
rect 10672 4483 10716 4491
rect 10258 4440 10273 4474
rect 10672 4466 10680 4483
rect 10697 4466 10716 4483
rect 10672 4458 10716 4466
rect 10294 4440 10309 4453
rect 10701 4440 10716 4458
rect 10737 4440 10752 4512
rect 10781 4440 10796 4564
rect 10825 4543 10840 4614
rect 11359 4597 11374 4614
rect 11349 4589 11382 4597
rect 11349 4572 11357 4589
rect 11374 4572 11382 4589
rect 11349 4564 11382 4572
rect 10817 4535 10850 4543
rect 10817 4518 10825 4535
rect 10842 4518 10850 4535
rect 10817 4510 10850 4518
rect 11250 4537 11283 4545
rect 11250 4520 11258 4537
rect 11275 4527 11283 4537
rect 11275 4520 11330 4527
rect 11250 4512 11330 4520
rect 10825 4440 10840 4510
rect 10916 4499 10949 4507
rect 10916 4489 10924 4499
rect 10869 4482 10924 4489
rect 10941 4482 10949 4499
rect 10869 4474 10949 4482
rect 11250 4483 11294 4491
rect 10869 4440 10884 4474
rect 11250 4466 11258 4483
rect 11275 4466 11294 4483
rect 11250 4458 11294 4466
rect 10905 4440 10920 4453
rect 11279 4440 11294 4458
rect 11315 4440 11330 4512
rect 11359 4440 11374 4564
rect 11403 4543 11418 4614
rect 11970 4597 11985 4614
rect 11960 4589 11993 4597
rect 11960 4572 11968 4589
rect 11985 4572 11993 4589
rect 11960 4564 11993 4572
rect 11395 4535 11428 4543
rect 11395 4518 11403 4535
rect 11420 4518 11428 4535
rect 11395 4510 11428 4518
rect 11861 4537 11894 4545
rect 11861 4520 11869 4537
rect 11886 4527 11894 4537
rect 11886 4520 11941 4527
rect 11861 4512 11941 4520
rect 11403 4440 11418 4510
rect 11494 4499 11527 4507
rect 11494 4489 11502 4499
rect 11447 4482 11502 4489
rect 11519 4482 11527 4499
rect 11447 4474 11527 4482
rect 11861 4483 11905 4491
rect 11447 4440 11462 4474
rect 11861 4466 11869 4483
rect 11886 4466 11905 4483
rect 11861 4458 11905 4466
rect 11483 4440 11498 4453
rect 11890 4440 11905 4458
rect 11926 4440 11941 4512
rect 11970 4440 11985 4564
rect 12014 4543 12029 4614
rect 12581 4597 12596 4614
rect 12571 4589 12604 4597
rect 12571 4572 12579 4589
rect 12596 4572 12604 4589
rect 12571 4564 12604 4572
rect 12006 4535 12039 4543
rect 12006 4518 12014 4535
rect 12031 4518 12039 4535
rect 12006 4510 12039 4518
rect 12472 4537 12505 4545
rect 12472 4520 12480 4537
rect 12497 4527 12505 4537
rect 12497 4520 12552 4527
rect 12472 4512 12552 4520
rect 12014 4440 12029 4510
rect 12105 4499 12138 4507
rect 12105 4489 12113 4499
rect 12058 4482 12113 4489
rect 12130 4482 12138 4499
rect 12058 4474 12138 4482
rect 12472 4483 12516 4491
rect 12058 4440 12073 4474
rect 12472 4466 12480 4483
rect 12497 4466 12516 4483
rect 12472 4458 12516 4466
rect 12094 4440 12109 4453
rect 12501 4440 12516 4458
rect 12537 4440 12552 4512
rect 12581 4440 12596 4564
rect 12625 4543 12640 4614
rect 12617 4535 12650 4543
rect 12617 4518 12625 4535
rect 12642 4518 12650 4535
rect 12617 4510 12650 4518
rect 12625 4440 12640 4510
rect 12716 4499 12749 4507
rect 12716 4489 12724 4499
rect 12669 4482 12724 4489
rect 12741 4482 12749 4499
rect 12669 4474 12749 4482
rect 12669 4440 12684 4474
rect 12705 4440 12720 4453
rect 9479 4306 9494 4340
rect 9515 4327 9530 4340
rect 9559 4327 9574 4340
rect 9603 4327 9618 4340
rect 9647 4327 9662 4340
rect 9683 4306 9698 4340
rect 9479 4291 9698 4306
rect 10090 4306 10105 4340
rect 10126 4327 10141 4340
rect 10170 4327 10185 4340
rect 10214 4327 10229 4340
rect 10258 4327 10273 4340
rect 10294 4306 10309 4340
rect 10090 4291 10309 4306
rect 10701 4306 10716 4340
rect 10737 4327 10752 4340
rect 10781 4327 10796 4340
rect 10825 4327 10840 4340
rect 10869 4327 10884 4340
rect 10905 4306 10920 4340
rect 10701 4291 10920 4306
rect 11279 4306 11294 4340
rect 11315 4327 11330 4340
rect 11359 4327 11374 4340
rect 11403 4327 11418 4340
rect 11447 4327 11462 4340
rect 11483 4306 11498 4340
rect 11279 4291 11498 4306
rect 11890 4306 11905 4340
rect 11926 4327 11941 4340
rect 11970 4327 11985 4340
rect 12014 4327 12029 4340
rect 12058 4327 12073 4340
rect 12094 4306 12109 4340
rect 11890 4291 12109 4306
rect 12501 4306 12516 4340
rect 12537 4327 12552 4340
rect 12581 4327 12596 4340
rect 12625 4327 12640 4340
rect 12669 4327 12684 4340
rect 12705 4306 12720 4340
rect 12501 4291 12720 4306
<< polycont >>
rect 10168 7802 10185 7819
rect 10069 7750 10086 7767
rect 10069 7696 10086 7713
rect 10779 7802 10796 7819
rect 10214 7748 10231 7765
rect 10680 7750 10697 7767
rect 10313 7712 10330 7729
rect 10680 7696 10697 7713
rect 11357 7802 11374 7819
rect 10825 7748 10842 7765
rect 11258 7750 11275 7767
rect 10924 7712 10941 7729
rect 11258 7696 11275 7713
rect 11968 7802 11985 7819
rect 11403 7748 11420 7765
rect 11869 7750 11886 7767
rect 11502 7712 11519 7729
rect 11869 7696 11886 7713
rect 12579 7802 12596 7819
rect 12014 7748 12031 7765
rect 12480 7750 12497 7767
rect 12113 7712 12130 7729
rect 12480 7696 12497 7713
rect 12625 7748 12642 7765
rect 12724 7712 12741 7729
rect 9557 7152 9574 7169
rect 9458 7100 9475 7117
rect 9458 7046 9475 7063
rect 10168 7152 10185 7169
rect 9603 7098 9620 7115
rect 10069 7100 10086 7117
rect 9702 7062 9719 7079
rect 10069 7046 10086 7063
rect 10779 7152 10796 7169
rect 10214 7098 10231 7115
rect 10680 7100 10697 7117
rect 10313 7062 10330 7079
rect 10680 7046 10697 7063
rect 11357 7152 11374 7169
rect 10825 7098 10842 7115
rect 11258 7100 11275 7117
rect 10924 7062 10941 7079
rect 11258 7046 11275 7063
rect 11968 7152 11985 7169
rect 11403 7098 11420 7115
rect 11869 7100 11886 7117
rect 11502 7062 11519 7079
rect 11869 7046 11886 7063
rect 12579 7152 12596 7169
rect 12014 7098 12031 7115
rect 12480 7100 12497 7117
rect 12113 7062 12130 7079
rect 12480 7046 12497 7063
rect 12625 7098 12642 7115
rect 12724 7062 12741 7079
rect 9557 6512 9574 6529
rect 9458 6460 9475 6477
rect 9458 6406 9475 6423
rect 10168 6512 10185 6529
rect 9603 6458 9620 6475
rect 10069 6460 10086 6477
rect 9702 6422 9719 6439
rect 10069 6406 10086 6423
rect 10779 6512 10796 6529
rect 10214 6458 10231 6475
rect 10680 6460 10697 6477
rect 10313 6422 10330 6439
rect 10680 6406 10697 6423
rect 11357 6512 11374 6529
rect 10825 6458 10842 6475
rect 11258 6460 11275 6477
rect 10924 6422 10941 6439
rect 11258 6406 11275 6423
rect 11968 6512 11985 6529
rect 11403 6458 11420 6475
rect 11869 6460 11886 6477
rect 11502 6422 11519 6439
rect 11869 6406 11886 6423
rect 12579 6512 12596 6529
rect 12014 6458 12031 6475
rect 12480 6460 12497 6477
rect 12113 6422 12130 6439
rect 12480 6406 12497 6423
rect 12625 6458 12642 6475
rect 12724 6422 12741 6439
rect 9557 5862 9574 5879
rect 9458 5810 9475 5827
rect 9458 5756 9475 5773
rect 10168 5862 10185 5879
rect 9603 5808 9620 5825
rect 10069 5810 10086 5827
rect 9702 5772 9719 5789
rect 10069 5756 10086 5773
rect 10779 5862 10796 5879
rect 10214 5808 10231 5825
rect 10680 5810 10697 5827
rect 10313 5772 10330 5789
rect 10680 5756 10697 5773
rect 11357 5862 11374 5879
rect 10825 5808 10842 5825
rect 11258 5810 11275 5827
rect 10924 5772 10941 5789
rect 11258 5756 11275 5773
rect 11968 5862 11985 5879
rect 11403 5808 11420 5825
rect 11869 5810 11886 5827
rect 11502 5772 11519 5789
rect 11869 5756 11886 5773
rect 12579 5862 12596 5879
rect 12014 5808 12031 5825
rect 12480 5810 12497 5827
rect 12113 5772 12130 5789
rect 12480 5756 12497 5773
rect 12625 5808 12642 5825
rect 12724 5772 12741 5789
rect 9557 5212 9574 5229
rect 9458 5160 9475 5177
rect 9458 5106 9475 5123
rect 10168 5212 10185 5229
rect 9603 5158 9620 5175
rect 10069 5160 10086 5177
rect 9702 5122 9719 5139
rect 10069 5106 10086 5123
rect 10779 5212 10796 5229
rect 10214 5158 10231 5175
rect 10680 5160 10697 5177
rect 10313 5122 10330 5139
rect 10680 5106 10697 5123
rect 11357 5212 11374 5229
rect 10825 5158 10842 5175
rect 11258 5160 11275 5177
rect 10924 5122 10941 5139
rect 11258 5106 11275 5123
rect 11968 5212 11985 5229
rect 11403 5158 11420 5175
rect 11869 5160 11886 5177
rect 11502 5122 11519 5139
rect 11869 5106 11886 5123
rect 12579 5212 12596 5229
rect 12014 5158 12031 5175
rect 12480 5160 12497 5177
rect 12113 5122 12130 5139
rect 12480 5106 12497 5123
rect 12625 5158 12642 5175
rect 12724 5122 12741 5139
rect 9557 4572 9574 4589
rect 9458 4520 9475 4537
rect 9458 4466 9475 4483
rect 10168 4572 10185 4589
rect 9603 4518 9620 4535
rect 10069 4520 10086 4537
rect 9702 4482 9719 4499
rect 10069 4466 10086 4483
rect 10779 4572 10796 4589
rect 10214 4518 10231 4535
rect 10680 4520 10697 4537
rect 10313 4482 10330 4499
rect 10680 4466 10697 4483
rect 11357 4572 11374 4589
rect 10825 4518 10842 4535
rect 11258 4520 11275 4537
rect 10924 4482 10941 4499
rect 11258 4466 11275 4483
rect 11968 4572 11985 4589
rect 11403 4518 11420 4535
rect 11869 4520 11886 4537
rect 11502 4482 11519 4499
rect 11869 4466 11886 4483
rect 12579 4572 12596 4589
rect 12014 4518 12031 4535
rect 12480 4520 12497 4537
rect 12113 4482 12130 4499
rect 12480 4466 12497 4483
rect 12625 4518 12642 4535
rect 12724 4482 12741 4499
<< locali >>
rect 10186 8062 10190 8081
rect 10209 8062 10213 8081
rect 10111 8039 10169 8047
rect 10111 8022 10147 8039
rect 10164 8022 10169 8039
rect 10111 8005 10169 8022
rect 10111 7988 10147 8005
rect 10164 7988 10169 8005
rect 10111 7971 10169 7988
rect 10111 7954 10147 7971
rect 10164 7954 10169 7971
rect 10111 7937 10169 7954
rect 10111 7920 10147 7937
rect 10164 7920 10169 7937
rect 10111 7903 10169 7920
rect 10111 7886 10147 7903
rect 10164 7886 10169 7903
rect 10111 7869 10169 7886
rect 10111 7852 10147 7869
rect 10164 7852 10169 7869
rect 10111 7844 10169 7852
rect 10186 8039 10213 8062
rect 10797 8062 10801 8081
rect 10820 8062 10824 8081
rect 10186 8022 10191 8039
rect 10208 8022 10213 8039
rect 10186 8005 10213 8022
rect 10186 7988 10191 8005
rect 10208 7988 10213 8005
rect 10186 7971 10213 7988
rect 10186 7954 10191 7971
rect 10208 7954 10213 7971
rect 10186 7937 10213 7954
rect 10186 7920 10191 7937
rect 10208 7920 10213 7937
rect 10186 7903 10213 7920
rect 10186 7886 10191 7903
rect 10208 7886 10213 7903
rect 10186 7869 10213 7886
rect 10186 7852 10191 7869
rect 10208 7852 10213 7869
rect 10186 7844 10213 7852
rect 10230 8039 10288 8047
rect 10230 8022 10235 8039
rect 10252 8022 10288 8039
rect 10230 8005 10288 8022
rect 10230 7988 10235 8005
rect 10252 7988 10288 8005
rect 10230 7971 10288 7988
rect 10230 7954 10235 7971
rect 10252 7954 10288 7971
rect 10230 7937 10288 7954
rect 10230 7920 10235 7937
rect 10252 7920 10288 7937
rect 10230 7903 10288 7920
rect 10230 7886 10235 7903
rect 10252 7886 10288 7903
rect 10230 7869 10288 7886
rect 10230 7852 10235 7869
rect 10252 7852 10288 7869
rect 10230 7844 10288 7852
rect 10061 7767 10094 7775
rect 10061 7750 10069 7767
rect 10086 7750 10094 7767
rect 10061 7742 10094 7750
rect 10111 7757 10138 7844
rect 10160 7819 10193 7827
rect 10160 7802 10168 7819
rect 10185 7811 10193 7819
rect 10261 7811 10288 7844
rect 10185 7802 10288 7811
rect 10160 7794 10288 7802
rect 10206 7765 10239 7773
rect 10206 7757 10214 7765
rect 10111 7748 10214 7757
rect 10231 7748 10239 7765
rect 10111 7740 10239 7748
rect 10061 7713 10094 7721
rect 10061 7696 10069 7713
rect 10086 7696 10094 7713
rect 10061 7688 10094 7696
rect 10111 7671 10138 7740
rect 10261 7671 10288 7794
rect 10722 8039 10780 8047
rect 10722 8022 10758 8039
rect 10775 8022 10780 8039
rect 10722 8005 10780 8022
rect 10722 7988 10758 8005
rect 10775 7988 10780 8005
rect 10722 7971 10780 7988
rect 10722 7954 10758 7971
rect 10775 7954 10780 7971
rect 10722 7937 10780 7954
rect 10722 7920 10758 7937
rect 10775 7920 10780 7937
rect 10722 7903 10780 7920
rect 10722 7886 10758 7903
rect 10775 7886 10780 7903
rect 10722 7869 10780 7886
rect 10722 7852 10758 7869
rect 10775 7852 10780 7869
rect 10722 7844 10780 7852
rect 10797 8039 10824 8062
rect 11375 8062 11379 8081
rect 11398 8062 11402 8081
rect 10797 8022 10802 8039
rect 10819 8022 10824 8039
rect 10797 8005 10824 8022
rect 10797 7988 10802 8005
rect 10819 7988 10824 8005
rect 10797 7971 10824 7988
rect 10797 7954 10802 7971
rect 10819 7954 10824 7971
rect 10797 7937 10824 7954
rect 10797 7920 10802 7937
rect 10819 7920 10824 7937
rect 10797 7903 10824 7920
rect 10797 7886 10802 7903
rect 10819 7886 10824 7903
rect 10797 7869 10824 7886
rect 10797 7852 10802 7869
rect 10819 7852 10824 7869
rect 10797 7844 10824 7852
rect 10841 8039 10899 8047
rect 10841 8022 10846 8039
rect 10863 8022 10899 8039
rect 10841 8005 10899 8022
rect 10841 7988 10846 8005
rect 10863 7988 10899 8005
rect 10841 7971 10899 7988
rect 10841 7954 10846 7971
rect 10863 7954 10899 7971
rect 10841 7937 10899 7954
rect 10841 7920 10846 7937
rect 10863 7920 10899 7937
rect 10841 7903 10899 7920
rect 10841 7886 10846 7903
rect 10863 7886 10899 7903
rect 10841 7869 10899 7886
rect 10841 7852 10846 7869
rect 10863 7852 10899 7869
rect 10841 7844 10899 7852
rect 10672 7767 10705 7775
rect 10672 7750 10680 7767
rect 10697 7750 10705 7767
rect 10672 7742 10705 7750
rect 10722 7757 10749 7844
rect 10771 7819 10804 7827
rect 10771 7802 10779 7819
rect 10796 7811 10804 7819
rect 10872 7811 10899 7844
rect 10796 7802 10899 7811
rect 10771 7794 10899 7802
rect 10817 7765 10850 7773
rect 10817 7757 10825 7765
rect 10722 7748 10825 7757
rect 10842 7748 10850 7765
rect 10722 7740 10850 7748
rect 10305 7729 10338 7737
rect 10305 7712 10313 7729
rect 10330 7712 10338 7729
rect 10305 7704 10338 7712
rect 10672 7713 10705 7721
rect 10672 7696 10680 7713
rect 10697 7696 10705 7713
rect 10672 7688 10705 7696
rect 10722 7671 10749 7740
rect 10872 7671 10899 7794
rect 11300 8039 11358 8047
rect 11300 8022 11336 8039
rect 11353 8022 11358 8039
rect 11300 8005 11358 8022
rect 11300 7988 11336 8005
rect 11353 7988 11358 8005
rect 11300 7971 11358 7988
rect 11300 7954 11336 7971
rect 11353 7954 11358 7971
rect 11300 7937 11358 7954
rect 11300 7920 11336 7937
rect 11353 7920 11358 7937
rect 11300 7903 11358 7920
rect 11300 7886 11336 7903
rect 11353 7886 11358 7903
rect 11300 7869 11358 7886
rect 11300 7852 11336 7869
rect 11353 7852 11358 7869
rect 11300 7844 11358 7852
rect 11375 8039 11402 8062
rect 11986 8062 11990 8081
rect 12009 8062 12013 8081
rect 11375 8022 11380 8039
rect 11397 8022 11402 8039
rect 11375 8005 11402 8022
rect 11375 7988 11380 8005
rect 11397 7988 11402 8005
rect 11375 7971 11402 7988
rect 11375 7954 11380 7971
rect 11397 7954 11402 7971
rect 11375 7937 11402 7954
rect 11375 7920 11380 7937
rect 11397 7920 11402 7937
rect 11375 7903 11402 7920
rect 11375 7886 11380 7903
rect 11397 7886 11402 7903
rect 11375 7869 11402 7886
rect 11375 7852 11380 7869
rect 11397 7852 11402 7869
rect 11375 7844 11402 7852
rect 11419 8039 11477 8047
rect 11419 8022 11424 8039
rect 11441 8022 11477 8039
rect 11419 8005 11477 8022
rect 11419 7988 11424 8005
rect 11441 7988 11477 8005
rect 11419 7971 11477 7988
rect 11419 7954 11424 7971
rect 11441 7954 11477 7971
rect 11419 7937 11477 7954
rect 11419 7920 11424 7937
rect 11441 7920 11477 7937
rect 11419 7903 11477 7920
rect 11419 7886 11424 7903
rect 11441 7886 11477 7903
rect 11419 7869 11477 7886
rect 11419 7852 11424 7869
rect 11441 7852 11477 7869
rect 11419 7844 11477 7852
rect 11250 7767 11283 7775
rect 11250 7750 11258 7767
rect 11275 7750 11283 7767
rect 11250 7742 11283 7750
rect 11300 7757 11327 7844
rect 11349 7819 11382 7827
rect 11349 7802 11357 7819
rect 11374 7811 11382 7819
rect 11450 7811 11477 7844
rect 11374 7802 11477 7811
rect 11349 7794 11477 7802
rect 11395 7765 11428 7773
rect 11395 7757 11403 7765
rect 11300 7748 11403 7757
rect 11420 7748 11428 7765
rect 11300 7740 11428 7748
rect 10916 7729 10949 7737
rect 10916 7712 10924 7729
rect 10941 7712 10949 7729
rect 10916 7704 10949 7712
rect 11250 7713 11283 7721
rect 11250 7696 11258 7713
rect 11275 7696 11283 7713
rect 11250 7688 11283 7696
rect 11300 7671 11327 7740
rect 11450 7671 11477 7794
rect 11911 8039 11969 8047
rect 11911 8022 11947 8039
rect 11964 8022 11969 8039
rect 11911 8005 11969 8022
rect 11911 7988 11947 8005
rect 11964 7988 11969 8005
rect 11911 7971 11969 7988
rect 11911 7954 11947 7971
rect 11964 7954 11969 7971
rect 11911 7937 11969 7954
rect 11911 7920 11947 7937
rect 11964 7920 11969 7937
rect 11911 7903 11969 7920
rect 11911 7886 11947 7903
rect 11964 7886 11969 7903
rect 11911 7869 11969 7886
rect 11911 7852 11947 7869
rect 11964 7852 11969 7869
rect 11911 7844 11969 7852
rect 11986 8039 12013 8062
rect 12597 8062 12601 8081
rect 12620 8062 12624 8081
rect 11986 8022 11991 8039
rect 12008 8022 12013 8039
rect 11986 8005 12013 8022
rect 11986 7988 11991 8005
rect 12008 7988 12013 8005
rect 11986 7971 12013 7988
rect 11986 7954 11991 7971
rect 12008 7954 12013 7971
rect 11986 7937 12013 7954
rect 11986 7920 11991 7937
rect 12008 7920 12013 7937
rect 11986 7903 12013 7920
rect 11986 7886 11991 7903
rect 12008 7886 12013 7903
rect 11986 7869 12013 7886
rect 11986 7852 11991 7869
rect 12008 7852 12013 7869
rect 11986 7844 12013 7852
rect 12030 8039 12088 8047
rect 12030 8022 12035 8039
rect 12052 8022 12088 8039
rect 12030 8005 12088 8022
rect 12030 7988 12035 8005
rect 12052 7988 12088 8005
rect 12030 7971 12088 7988
rect 12030 7954 12035 7971
rect 12052 7954 12088 7971
rect 12030 7937 12088 7954
rect 12030 7920 12035 7937
rect 12052 7920 12088 7937
rect 12030 7903 12088 7920
rect 12030 7886 12035 7903
rect 12052 7886 12088 7903
rect 12030 7869 12088 7886
rect 12030 7852 12035 7869
rect 12052 7852 12088 7869
rect 12030 7844 12088 7852
rect 11861 7767 11894 7775
rect 11861 7750 11869 7767
rect 11886 7750 11894 7767
rect 11861 7742 11894 7750
rect 11911 7757 11938 7844
rect 11960 7819 11993 7827
rect 11960 7802 11968 7819
rect 11985 7811 11993 7819
rect 12061 7811 12088 7844
rect 11985 7802 12088 7811
rect 11960 7794 12088 7802
rect 12006 7765 12039 7773
rect 12006 7757 12014 7765
rect 11911 7748 12014 7757
rect 12031 7748 12039 7765
rect 11911 7740 12039 7748
rect 11494 7729 11527 7737
rect 11494 7712 11502 7729
rect 11519 7712 11527 7729
rect 11494 7704 11527 7712
rect 11861 7713 11894 7721
rect 11861 7696 11869 7713
rect 11886 7696 11894 7713
rect 11861 7688 11894 7696
rect 11911 7671 11938 7740
rect 12061 7671 12088 7794
rect 12522 8039 12580 8047
rect 12522 8022 12558 8039
rect 12575 8022 12580 8039
rect 12522 8005 12580 8022
rect 12522 7988 12558 8005
rect 12575 7988 12580 8005
rect 12522 7971 12580 7988
rect 12522 7954 12558 7971
rect 12575 7954 12580 7971
rect 12522 7937 12580 7954
rect 12522 7920 12558 7937
rect 12575 7920 12580 7937
rect 12522 7903 12580 7920
rect 12522 7886 12558 7903
rect 12575 7886 12580 7903
rect 12522 7869 12580 7886
rect 12522 7852 12558 7869
rect 12575 7852 12580 7869
rect 12522 7844 12580 7852
rect 12597 8039 12624 8062
rect 12597 8022 12602 8039
rect 12619 8022 12624 8039
rect 12597 8005 12624 8022
rect 12597 7988 12602 8005
rect 12619 7988 12624 8005
rect 12597 7971 12624 7988
rect 12597 7954 12602 7971
rect 12619 7954 12624 7971
rect 12597 7937 12624 7954
rect 12597 7920 12602 7937
rect 12619 7920 12624 7937
rect 12597 7903 12624 7920
rect 12597 7886 12602 7903
rect 12619 7886 12624 7903
rect 12597 7869 12624 7886
rect 12597 7852 12602 7869
rect 12619 7852 12624 7869
rect 12597 7844 12624 7852
rect 12641 8039 12699 8047
rect 12641 8022 12646 8039
rect 12663 8022 12699 8039
rect 12641 8005 12699 8022
rect 12641 7988 12646 8005
rect 12663 7988 12699 8005
rect 12641 7971 12699 7988
rect 12641 7954 12646 7971
rect 12663 7954 12699 7971
rect 12641 7937 12699 7954
rect 12641 7920 12646 7937
rect 12663 7920 12699 7937
rect 12641 7903 12699 7920
rect 12641 7886 12646 7903
rect 12663 7886 12699 7903
rect 12641 7869 12699 7886
rect 12641 7852 12646 7869
rect 12663 7852 12699 7869
rect 12641 7844 12699 7852
rect 12472 7767 12505 7775
rect 12472 7750 12480 7767
rect 12497 7750 12505 7767
rect 12472 7742 12505 7750
rect 12522 7757 12549 7844
rect 12571 7819 12604 7827
rect 12571 7802 12579 7819
rect 12596 7811 12604 7819
rect 12672 7811 12699 7844
rect 12596 7802 12699 7811
rect 12571 7794 12699 7802
rect 12617 7765 12650 7773
rect 12617 7757 12625 7765
rect 12522 7748 12625 7757
rect 12642 7748 12650 7765
rect 12522 7740 12650 7748
rect 12105 7729 12138 7737
rect 12105 7712 12113 7729
rect 12130 7712 12138 7729
rect 12105 7704 12138 7712
rect 12472 7713 12505 7721
rect 12472 7696 12480 7713
rect 12497 7696 12505 7713
rect 12472 7688 12505 7696
rect 12522 7671 12549 7740
rect 12672 7671 12699 7794
rect 12716 7729 12749 7737
rect 12716 7712 12724 7729
rect 12741 7712 12749 7729
rect 12716 7704 12749 7712
rect 10062 7663 10089 7671
rect 10062 7646 10067 7663
rect 10084 7646 10089 7663
rect 10062 7629 10089 7646
rect 10062 7612 10067 7629
rect 10084 7612 10089 7629
rect 10062 7595 10089 7612
rect 10062 7578 10067 7595
rect 10084 7578 10089 7595
rect 10062 7570 10089 7578
rect 10111 7663 10169 7671
rect 10111 7646 10147 7663
rect 10164 7646 10169 7663
rect 10111 7629 10169 7646
rect 10111 7612 10147 7629
rect 10164 7612 10169 7629
rect 10111 7595 10169 7612
rect 10111 7578 10147 7595
rect 10164 7578 10169 7595
rect 10111 7570 10169 7578
rect 10186 7663 10213 7671
rect 10186 7646 10191 7663
rect 10208 7646 10213 7663
rect 10186 7629 10213 7646
rect 10186 7612 10191 7629
rect 10208 7612 10213 7629
rect 10186 7595 10213 7612
rect 10186 7578 10191 7595
rect 10208 7578 10213 7595
rect 10186 7555 10213 7578
rect 10230 7663 10288 7671
rect 10230 7646 10235 7663
rect 10252 7646 10288 7663
rect 10230 7629 10288 7646
rect 10230 7612 10235 7629
rect 10252 7612 10288 7629
rect 10230 7595 10288 7612
rect 10230 7578 10235 7595
rect 10252 7578 10288 7595
rect 10230 7570 10288 7578
rect 10310 7663 10337 7671
rect 10310 7646 10315 7663
rect 10332 7646 10337 7663
rect 10310 7629 10337 7646
rect 10310 7612 10315 7629
rect 10332 7612 10337 7629
rect 10310 7595 10337 7612
rect 10310 7578 10315 7595
rect 10332 7578 10337 7595
rect 10310 7570 10337 7578
rect 10673 7663 10700 7671
rect 10673 7646 10678 7663
rect 10695 7646 10700 7663
rect 10673 7629 10700 7646
rect 10673 7612 10678 7629
rect 10695 7612 10700 7629
rect 10673 7595 10700 7612
rect 10673 7578 10678 7595
rect 10695 7578 10700 7595
rect 10673 7570 10700 7578
rect 10722 7663 10780 7671
rect 10722 7646 10758 7663
rect 10775 7646 10780 7663
rect 10722 7629 10780 7646
rect 10722 7612 10758 7629
rect 10775 7612 10780 7629
rect 10722 7595 10780 7612
rect 10722 7578 10758 7595
rect 10775 7578 10780 7595
rect 10722 7570 10780 7578
rect 10797 7663 10824 7671
rect 10797 7646 10802 7663
rect 10819 7646 10824 7663
rect 10797 7629 10824 7646
rect 10797 7612 10802 7629
rect 10819 7612 10824 7629
rect 10797 7595 10824 7612
rect 10797 7578 10802 7595
rect 10819 7578 10824 7595
rect 10186 7536 10190 7555
rect 10209 7536 10213 7555
rect 10797 7555 10824 7578
rect 10841 7663 10899 7671
rect 10841 7646 10846 7663
rect 10863 7646 10899 7663
rect 10841 7629 10899 7646
rect 10841 7612 10846 7629
rect 10863 7612 10899 7629
rect 10841 7595 10899 7612
rect 10841 7578 10846 7595
rect 10863 7578 10899 7595
rect 10841 7570 10899 7578
rect 10921 7663 10948 7671
rect 10921 7646 10926 7663
rect 10943 7646 10948 7663
rect 10921 7629 10948 7646
rect 10921 7612 10926 7629
rect 10943 7612 10948 7629
rect 10921 7595 10948 7612
rect 10921 7578 10926 7595
rect 10943 7578 10948 7595
rect 10921 7570 10948 7578
rect 11251 7663 11278 7671
rect 11251 7646 11256 7663
rect 11273 7646 11278 7663
rect 11251 7629 11278 7646
rect 11251 7612 11256 7629
rect 11273 7612 11278 7629
rect 11251 7595 11278 7612
rect 11251 7578 11256 7595
rect 11273 7578 11278 7595
rect 11251 7570 11278 7578
rect 11300 7663 11358 7671
rect 11300 7646 11336 7663
rect 11353 7646 11358 7663
rect 11300 7629 11358 7646
rect 11300 7612 11336 7629
rect 11353 7612 11358 7629
rect 11300 7595 11358 7612
rect 11300 7578 11336 7595
rect 11353 7578 11358 7595
rect 11300 7570 11358 7578
rect 11375 7663 11402 7671
rect 11375 7646 11380 7663
rect 11397 7646 11402 7663
rect 11375 7629 11402 7646
rect 11375 7612 11380 7629
rect 11397 7612 11402 7629
rect 11375 7595 11402 7612
rect 11375 7578 11380 7595
rect 11397 7578 11402 7595
rect 10797 7536 10801 7555
rect 10820 7536 10824 7555
rect 11375 7555 11402 7578
rect 11419 7663 11477 7671
rect 11419 7646 11424 7663
rect 11441 7646 11477 7663
rect 11419 7629 11477 7646
rect 11419 7612 11424 7629
rect 11441 7612 11477 7629
rect 11419 7595 11477 7612
rect 11419 7578 11424 7595
rect 11441 7578 11477 7595
rect 11419 7570 11477 7578
rect 11499 7663 11526 7671
rect 11499 7646 11504 7663
rect 11521 7646 11526 7663
rect 11499 7629 11526 7646
rect 11499 7612 11504 7629
rect 11521 7612 11526 7629
rect 11499 7595 11526 7612
rect 11499 7578 11504 7595
rect 11521 7578 11526 7595
rect 11499 7570 11526 7578
rect 11862 7663 11889 7671
rect 11862 7646 11867 7663
rect 11884 7646 11889 7663
rect 11862 7629 11889 7646
rect 11862 7612 11867 7629
rect 11884 7612 11889 7629
rect 11862 7595 11889 7612
rect 11862 7578 11867 7595
rect 11884 7578 11889 7595
rect 11862 7570 11889 7578
rect 11911 7663 11969 7671
rect 11911 7646 11947 7663
rect 11964 7646 11969 7663
rect 11911 7629 11969 7646
rect 11911 7612 11947 7629
rect 11964 7612 11969 7629
rect 11911 7595 11969 7612
rect 11911 7578 11947 7595
rect 11964 7578 11969 7595
rect 11911 7570 11969 7578
rect 11986 7663 12013 7671
rect 11986 7646 11991 7663
rect 12008 7646 12013 7663
rect 11986 7629 12013 7646
rect 11986 7612 11991 7629
rect 12008 7612 12013 7629
rect 11986 7595 12013 7612
rect 11986 7578 11991 7595
rect 12008 7578 12013 7595
rect 11375 7536 11379 7555
rect 11398 7536 11402 7555
rect 11986 7555 12013 7578
rect 12030 7663 12088 7671
rect 12030 7646 12035 7663
rect 12052 7646 12088 7663
rect 12030 7629 12088 7646
rect 12030 7612 12035 7629
rect 12052 7612 12088 7629
rect 12030 7595 12088 7612
rect 12030 7578 12035 7595
rect 12052 7578 12088 7595
rect 12030 7570 12088 7578
rect 12110 7663 12137 7671
rect 12110 7646 12115 7663
rect 12132 7646 12137 7663
rect 12110 7629 12137 7646
rect 12110 7612 12115 7629
rect 12132 7612 12137 7629
rect 12110 7595 12137 7612
rect 12110 7578 12115 7595
rect 12132 7578 12137 7595
rect 12110 7570 12137 7578
rect 12473 7663 12500 7671
rect 12473 7646 12478 7663
rect 12495 7646 12500 7663
rect 12473 7629 12500 7646
rect 12473 7612 12478 7629
rect 12495 7612 12500 7629
rect 12473 7595 12500 7612
rect 12473 7578 12478 7595
rect 12495 7578 12500 7595
rect 12473 7570 12500 7578
rect 12522 7663 12580 7671
rect 12522 7646 12558 7663
rect 12575 7646 12580 7663
rect 12522 7629 12580 7646
rect 12522 7612 12558 7629
rect 12575 7612 12580 7629
rect 12522 7595 12580 7612
rect 12522 7578 12558 7595
rect 12575 7578 12580 7595
rect 12522 7570 12580 7578
rect 12597 7663 12624 7671
rect 12597 7646 12602 7663
rect 12619 7646 12624 7663
rect 12597 7629 12624 7646
rect 12597 7612 12602 7629
rect 12619 7612 12624 7629
rect 12597 7595 12624 7612
rect 12597 7578 12602 7595
rect 12619 7578 12624 7595
rect 11986 7536 11990 7555
rect 12009 7536 12013 7555
rect 12597 7555 12624 7578
rect 12641 7663 12699 7671
rect 12641 7646 12646 7663
rect 12663 7646 12699 7663
rect 12641 7629 12699 7646
rect 12641 7612 12646 7629
rect 12663 7612 12699 7629
rect 12641 7595 12699 7612
rect 12641 7578 12646 7595
rect 12663 7578 12699 7595
rect 12641 7570 12699 7578
rect 12721 7663 12748 7671
rect 12721 7646 12726 7663
rect 12743 7646 12748 7663
rect 12721 7629 12748 7646
rect 12721 7612 12726 7629
rect 12743 7612 12748 7629
rect 12721 7595 12748 7612
rect 12721 7578 12726 7595
rect 12743 7578 12748 7595
rect 12721 7570 12748 7578
rect 12597 7536 12601 7555
rect 12620 7536 12624 7555
rect 9575 7412 9579 7431
rect 9598 7412 9602 7431
rect 9500 7389 9558 7397
rect 9500 7372 9536 7389
rect 9553 7372 9558 7389
rect 9500 7355 9558 7372
rect 9500 7338 9536 7355
rect 9553 7338 9558 7355
rect 9500 7321 9558 7338
rect 9500 7304 9536 7321
rect 9553 7304 9558 7321
rect 9500 7287 9558 7304
rect 9500 7270 9536 7287
rect 9553 7270 9558 7287
rect 9500 7253 9558 7270
rect 9500 7236 9536 7253
rect 9553 7236 9558 7253
rect 9500 7219 9558 7236
rect 9500 7202 9536 7219
rect 9553 7202 9558 7219
rect 9500 7194 9558 7202
rect 9575 7389 9602 7412
rect 10186 7412 10190 7431
rect 10209 7412 10213 7431
rect 9575 7372 9580 7389
rect 9597 7372 9602 7389
rect 9575 7355 9602 7372
rect 9575 7338 9580 7355
rect 9597 7338 9602 7355
rect 9575 7321 9602 7338
rect 9575 7304 9580 7321
rect 9597 7304 9602 7321
rect 9575 7287 9602 7304
rect 9575 7270 9580 7287
rect 9597 7270 9602 7287
rect 9575 7253 9602 7270
rect 9575 7236 9580 7253
rect 9597 7236 9602 7253
rect 9575 7219 9602 7236
rect 9575 7202 9580 7219
rect 9597 7202 9602 7219
rect 9575 7194 9602 7202
rect 9619 7389 9677 7397
rect 9619 7372 9624 7389
rect 9641 7372 9677 7389
rect 9619 7355 9677 7372
rect 9619 7338 9624 7355
rect 9641 7338 9677 7355
rect 9619 7321 9677 7338
rect 9619 7304 9624 7321
rect 9641 7304 9677 7321
rect 9619 7287 9677 7304
rect 9619 7270 9624 7287
rect 9641 7270 9677 7287
rect 9619 7253 9677 7270
rect 9619 7236 9624 7253
rect 9641 7236 9677 7253
rect 9619 7219 9677 7236
rect 9619 7202 9624 7219
rect 9641 7202 9677 7219
rect 9619 7194 9677 7202
rect 9450 7117 9483 7125
rect 9450 7100 9458 7117
rect 9475 7100 9483 7117
rect 9450 7092 9483 7100
rect 9500 7107 9527 7194
rect 9549 7169 9582 7177
rect 9549 7152 9557 7169
rect 9574 7161 9582 7169
rect 9650 7161 9677 7194
rect 9574 7152 9677 7161
rect 9549 7144 9677 7152
rect 9595 7115 9628 7123
rect 9595 7107 9603 7115
rect 9500 7098 9603 7107
rect 9620 7098 9628 7115
rect 9500 7090 9628 7098
rect 9450 7063 9483 7071
rect 9450 7046 9458 7063
rect 9475 7046 9483 7063
rect 9450 7038 9483 7046
rect 9500 7021 9527 7090
rect 9650 7021 9677 7144
rect 10111 7389 10169 7397
rect 10111 7372 10147 7389
rect 10164 7372 10169 7389
rect 10111 7355 10169 7372
rect 10111 7338 10147 7355
rect 10164 7338 10169 7355
rect 10111 7321 10169 7338
rect 10111 7304 10147 7321
rect 10164 7304 10169 7321
rect 10111 7287 10169 7304
rect 10111 7270 10147 7287
rect 10164 7270 10169 7287
rect 10111 7253 10169 7270
rect 10111 7236 10147 7253
rect 10164 7236 10169 7253
rect 10111 7219 10169 7236
rect 10111 7202 10147 7219
rect 10164 7202 10169 7219
rect 10111 7194 10169 7202
rect 10186 7389 10213 7412
rect 10797 7412 10801 7431
rect 10820 7412 10824 7431
rect 10186 7372 10191 7389
rect 10208 7372 10213 7389
rect 10186 7355 10213 7372
rect 10186 7338 10191 7355
rect 10208 7338 10213 7355
rect 10186 7321 10213 7338
rect 10186 7304 10191 7321
rect 10208 7304 10213 7321
rect 10186 7287 10213 7304
rect 10186 7270 10191 7287
rect 10208 7270 10213 7287
rect 10186 7253 10213 7270
rect 10186 7236 10191 7253
rect 10208 7236 10213 7253
rect 10186 7219 10213 7236
rect 10186 7202 10191 7219
rect 10208 7202 10213 7219
rect 10186 7194 10213 7202
rect 10230 7389 10288 7397
rect 10230 7372 10235 7389
rect 10252 7372 10288 7389
rect 10230 7355 10288 7372
rect 10230 7338 10235 7355
rect 10252 7338 10288 7355
rect 10230 7321 10288 7338
rect 10230 7304 10235 7321
rect 10252 7304 10288 7321
rect 10230 7287 10288 7304
rect 10230 7270 10235 7287
rect 10252 7270 10288 7287
rect 10230 7253 10288 7270
rect 10230 7236 10235 7253
rect 10252 7236 10288 7253
rect 10230 7219 10288 7236
rect 10230 7202 10235 7219
rect 10252 7202 10288 7219
rect 10230 7194 10288 7202
rect 10061 7117 10094 7125
rect 10061 7100 10069 7117
rect 10086 7100 10094 7117
rect 10061 7092 10094 7100
rect 10111 7107 10138 7194
rect 10160 7169 10193 7177
rect 10160 7152 10168 7169
rect 10185 7161 10193 7169
rect 10261 7161 10288 7194
rect 10185 7152 10288 7161
rect 10160 7144 10288 7152
rect 10206 7115 10239 7123
rect 10206 7107 10214 7115
rect 10111 7098 10214 7107
rect 10231 7098 10239 7115
rect 10111 7090 10239 7098
rect 9694 7079 9727 7087
rect 9694 7062 9702 7079
rect 9719 7062 9727 7079
rect 9694 7054 9727 7062
rect 10061 7063 10094 7071
rect 10061 7046 10069 7063
rect 10086 7046 10094 7063
rect 10061 7038 10094 7046
rect 10111 7021 10138 7090
rect 10261 7021 10288 7144
rect 10722 7389 10780 7397
rect 10722 7372 10758 7389
rect 10775 7372 10780 7389
rect 10722 7355 10780 7372
rect 10722 7338 10758 7355
rect 10775 7338 10780 7355
rect 10722 7321 10780 7338
rect 10722 7304 10758 7321
rect 10775 7304 10780 7321
rect 10722 7287 10780 7304
rect 10722 7270 10758 7287
rect 10775 7270 10780 7287
rect 10722 7253 10780 7270
rect 10722 7236 10758 7253
rect 10775 7236 10780 7253
rect 10722 7219 10780 7236
rect 10722 7202 10758 7219
rect 10775 7202 10780 7219
rect 10722 7194 10780 7202
rect 10797 7389 10824 7412
rect 11375 7412 11379 7431
rect 11398 7412 11402 7431
rect 10797 7372 10802 7389
rect 10819 7372 10824 7389
rect 10797 7355 10824 7372
rect 10797 7338 10802 7355
rect 10819 7338 10824 7355
rect 10797 7321 10824 7338
rect 10797 7304 10802 7321
rect 10819 7304 10824 7321
rect 10797 7287 10824 7304
rect 10797 7270 10802 7287
rect 10819 7270 10824 7287
rect 10797 7253 10824 7270
rect 10797 7236 10802 7253
rect 10819 7236 10824 7253
rect 10797 7219 10824 7236
rect 10797 7202 10802 7219
rect 10819 7202 10824 7219
rect 10797 7194 10824 7202
rect 10841 7389 10899 7397
rect 10841 7372 10846 7389
rect 10863 7372 10899 7389
rect 10841 7355 10899 7372
rect 10841 7338 10846 7355
rect 10863 7338 10899 7355
rect 10841 7321 10899 7338
rect 10841 7304 10846 7321
rect 10863 7304 10899 7321
rect 10841 7287 10899 7304
rect 10841 7270 10846 7287
rect 10863 7270 10899 7287
rect 10841 7253 10899 7270
rect 10841 7236 10846 7253
rect 10863 7236 10899 7253
rect 10841 7219 10899 7236
rect 10841 7202 10846 7219
rect 10863 7202 10899 7219
rect 10841 7194 10899 7202
rect 10672 7117 10705 7125
rect 10672 7100 10680 7117
rect 10697 7100 10705 7117
rect 10672 7092 10705 7100
rect 10722 7107 10749 7194
rect 10771 7169 10804 7177
rect 10771 7152 10779 7169
rect 10796 7161 10804 7169
rect 10872 7161 10899 7194
rect 10796 7152 10899 7161
rect 10771 7144 10899 7152
rect 10817 7115 10850 7123
rect 10817 7107 10825 7115
rect 10722 7098 10825 7107
rect 10842 7098 10850 7115
rect 10722 7090 10850 7098
rect 10305 7079 10338 7087
rect 10305 7062 10313 7079
rect 10330 7062 10338 7079
rect 10305 7054 10338 7062
rect 10672 7063 10705 7071
rect 10672 7046 10680 7063
rect 10697 7046 10705 7063
rect 10672 7038 10705 7046
rect 10722 7021 10749 7090
rect 10872 7021 10899 7144
rect 11300 7389 11358 7397
rect 11300 7372 11336 7389
rect 11353 7372 11358 7389
rect 11300 7355 11358 7372
rect 11300 7338 11336 7355
rect 11353 7338 11358 7355
rect 11300 7321 11358 7338
rect 11300 7304 11336 7321
rect 11353 7304 11358 7321
rect 11300 7287 11358 7304
rect 11300 7270 11336 7287
rect 11353 7270 11358 7287
rect 11300 7253 11358 7270
rect 11300 7236 11336 7253
rect 11353 7236 11358 7253
rect 11300 7219 11358 7236
rect 11300 7202 11336 7219
rect 11353 7202 11358 7219
rect 11300 7194 11358 7202
rect 11375 7389 11402 7412
rect 11986 7412 11990 7431
rect 12009 7412 12013 7431
rect 11375 7372 11380 7389
rect 11397 7372 11402 7389
rect 11375 7355 11402 7372
rect 11375 7338 11380 7355
rect 11397 7338 11402 7355
rect 11375 7321 11402 7338
rect 11375 7304 11380 7321
rect 11397 7304 11402 7321
rect 11375 7287 11402 7304
rect 11375 7270 11380 7287
rect 11397 7270 11402 7287
rect 11375 7253 11402 7270
rect 11375 7236 11380 7253
rect 11397 7236 11402 7253
rect 11375 7219 11402 7236
rect 11375 7202 11380 7219
rect 11397 7202 11402 7219
rect 11375 7194 11402 7202
rect 11419 7389 11477 7397
rect 11419 7372 11424 7389
rect 11441 7372 11477 7389
rect 11419 7355 11477 7372
rect 11419 7338 11424 7355
rect 11441 7338 11477 7355
rect 11419 7321 11477 7338
rect 11419 7304 11424 7321
rect 11441 7304 11477 7321
rect 11419 7287 11477 7304
rect 11419 7270 11424 7287
rect 11441 7270 11477 7287
rect 11419 7253 11477 7270
rect 11419 7236 11424 7253
rect 11441 7236 11477 7253
rect 11419 7219 11477 7236
rect 11419 7202 11424 7219
rect 11441 7202 11477 7219
rect 11419 7194 11477 7202
rect 11250 7117 11283 7125
rect 11250 7100 11258 7117
rect 11275 7100 11283 7117
rect 11250 7092 11283 7100
rect 11300 7107 11327 7194
rect 11349 7169 11382 7177
rect 11349 7152 11357 7169
rect 11374 7161 11382 7169
rect 11450 7161 11477 7194
rect 11374 7152 11477 7161
rect 11349 7144 11477 7152
rect 11395 7115 11428 7123
rect 11395 7107 11403 7115
rect 11300 7098 11403 7107
rect 11420 7098 11428 7115
rect 11300 7090 11428 7098
rect 10916 7079 10949 7087
rect 10916 7062 10924 7079
rect 10941 7062 10949 7079
rect 10916 7054 10949 7062
rect 11250 7063 11283 7071
rect 11250 7046 11258 7063
rect 11275 7046 11283 7063
rect 11250 7038 11283 7046
rect 11300 7021 11327 7090
rect 11450 7021 11477 7144
rect 11911 7389 11969 7397
rect 11911 7372 11947 7389
rect 11964 7372 11969 7389
rect 11911 7355 11969 7372
rect 11911 7338 11947 7355
rect 11964 7338 11969 7355
rect 11911 7321 11969 7338
rect 11911 7304 11947 7321
rect 11964 7304 11969 7321
rect 11911 7287 11969 7304
rect 11911 7270 11947 7287
rect 11964 7270 11969 7287
rect 11911 7253 11969 7270
rect 11911 7236 11947 7253
rect 11964 7236 11969 7253
rect 11911 7219 11969 7236
rect 11911 7202 11947 7219
rect 11964 7202 11969 7219
rect 11911 7194 11969 7202
rect 11986 7389 12013 7412
rect 12597 7412 12601 7431
rect 12620 7412 12624 7431
rect 11986 7372 11991 7389
rect 12008 7372 12013 7389
rect 11986 7355 12013 7372
rect 11986 7338 11991 7355
rect 12008 7338 12013 7355
rect 11986 7321 12013 7338
rect 11986 7304 11991 7321
rect 12008 7304 12013 7321
rect 11986 7287 12013 7304
rect 11986 7270 11991 7287
rect 12008 7270 12013 7287
rect 11986 7253 12013 7270
rect 11986 7236 11991 7253
rect 12008 7236 12013 7253
rect 11986 7219 12013 7236
rect 11986 7202 11991 7219
rect 12008 7202 12013 7219
rect 11986 7194 12013 7202
rect 12030 7389 12088 7397
rect 12030 7372 12035 7389
rect 12052 7372 12088 7389
rect 12030 7355 12088 7372
rect 12030 7338 12035 7355
rect 12052 7338 12088 7355
rect 12030 7321 12088 7338
rect 12030 7304 12035 7321
rect 12052 7304 12088 7321
rect 12030 7287 12088 7304
rect 12030 7270 12035 7287
rect 12052 7270 12088 7287
rect 12030 7253 12088 7270
rect 12030 7236 12035 7253
rect 12052 7236 12088 7253
rect 12030 7219 12088 7236
rect 12030 7202 12035 7219
rect 12052 7202 12088 7219
rect 12030 7194 12088 7202
rect 11861 7117 11894 7125
rect 11861 7100 11869 7117
rect 11886 7100 11894 7117
rect 11861 7092 11894 7100
rect 11911 7107 11938 7194
rect 11960 7169 11993 7177
rect 11960 7152 11968 7169
rect 11985 7161 11993 7169
rect 12061 7161 12088 7194
rect 11985 7152 12088 7161
rect 11960 7144 12088 7152
rect 12006 7115 12039 7123
rect 12006 7107 12014 7115
rect 11911 7098 12014 7107
rect 12031 7098 12039 7115
rect 11911 7090 12039 7098
rect 11494 7079 11527 7087
rect 11494 7062 11502 7079
rect 11519 7062 11527 7079
rect 11494 7054 11527 7062
rect 11861 7063 11894 7071
rect 11861 7046 11869 7063
rect 11886 7046 11894 7063
rect 11861 7038 11894 7046
rect 11911 7021 11938 7090
rect 12061 7021 12088 7144
rect 12522 7389 12580 7397
rect 12522 7372 12558 7389
rect 12575 7372 12580 7389
rect 12522 7355 12580 7372
rect 12522 7338 12558 7355
rect 12575 7338 12580 7355
rect 12522 7321 12580 7338
rect 12522 7304 12558 7321
rect 12575 7304 12580 7321
rect 12522 7287 12580 7304
rect 12522 7270 12558 7287
rect 12575 7270 12580 7287
rect 12522 7253 12580 7270
rect 12522 7236 12558 7253
rect 12575 7236 12580 7253
rect 12522 7219 12580 7236
rect 12522 7202 12558 7219
rect 12575 7202 12580 7219
rect 12522 7194 12580 7202
rect 12597 7389 12624 7412
rect 12597 7372 12602 7389
rect 12619 7372 12624 7389
rect 12597 7355 12624 7372
rect 12597 7338 12602 7355
rect 12619 7338 12624 7355
rect 12597 7321 12624 7338
rect 12597 7304 12602 7321
rect 12619 7304 12624 7321
rect 12597 7287 12624 7304
rect 12597 7270 12602 7287
rect 12619 7270 12624 7287
rect 12597 7253 12624 7270
rect 12597 7236 12602 7253
rect 12619 7236 12624 7253
rect 12597 7219 12624 7236
rect 12597 7202 12602 7219
rect 12619 7202 12624 7219
rect 12597 7194 12624 7202
rect 12641 7389 12699 7397
rect 12641 7372 12646 7389
rect 12663 7372 12699 7389
rect 12641 7355 12699 7372
rect 12641 7338 12646 7355
rect 12663 7338 12699 7355
rect 12641 7321 12699 7338
rect 12641 7304 12646 7321
rect 12663 7304 12699 7321
rect 12641 7287 12699 7304
rect 12641 7270 12646 7287
rect 12663 7270 12699 7287
rect 12641 7253 12699 7270
rect 12641 7236 12646 7253
rect 12663 7236 12699 7253
rect 12641 7219 12699 7236
rect 12641 7202 12646 7219
rect 12663 7202 12699 7219
rect 12641 7194 12699 7202
rect 12472 7117 12505 7125
rect 12472 7100 12480 7117
rect 12497 7100 12505 7117
rect 12472 7092 12505 7100
rect 12522 7107 12549 7194
rect 12571 7169 12604 7177
rect 12571 7152 12579 7169
rect 12596 7161 12604 7169
rect 12672 7161 12699 7194
rect 12596 7152 12699 7161
rect 12571 7144 12699 7152
rect 12617 7115 12650 7123
rect 12617 7107 12625 7115
rect 12522 7098 12625 7107
rect 12642 7098 12650 7115
rect 12522 7090 12650 7098
rect 12105 7079 12138 7087
rect 12105 7062 12113 7079
rect 12130 7062 12138 7079
rect 12105 7054 12138 7062
rect 12472 7063 12505 7071
rect 12472 7046 12480 7063
rect 12497 7046 12505 7063
rect 12472 7038 12505 7046
rect 12522 7021 12549 7090
rect 12672 7021 12699 7144
rect 12716 7079 12749 7087
rect 12716 7062 12724 7079
rect 12741 7062 12749 7079
rect 12716 7054 12749 7062
rect 9451 7013 9478 7021
rect 9451 6996 9456 7013
rect 9473 6996 9478 7013
rect 9451 6979 9478 6996
rect 9451 6962 9456 6979
rect 9473 6962 9478 6979
rect 9451 6945 9478 6962
rect 9451 6928 9456 6945
rect 9473 6928 9478 6945
rect 9451 6920 9478 6928
rect 9500 7013 9558 7021
rect 9500 6996 9536 7013
rect 9553 6996 9558 7013
rect 9500 6979 9558 6996
rect 9500 6962 9536 6979
rect 9553 6962 9558 6979
rect 9500 6945 9558 6962
rect 9500 6928 9536 6945
rect 9553 6928 9558 6945
rect 9500 6920 9558 6928
rect 9575 7013 9602 7021
rect 9575 6996 9580 7013
rect 9597 6996 9602 7013
rect 9575 6979 9602 6996
rect 9575 6962 9580 6979
rect 9597 6962 9602 6979
rect 9575 6945 9602 6962
rect 9575 6928 9580 6945
rect 9597 6928 9602 6945
rect 9575 6905 9602 6928
rect 9619 7013 9677 7021
rect 9619 6996 9624 7013
rect 9641 6996 9677 7013
rect 9619 6979 9677 6996
rect 9619 6962 9624 6979
rect 9641 6962 9677 6979
rect 9619 6945 9677 6962
rect 9619 6928 9624 6945
rect 9641 6928 9677 6945
rect 9619 6920 9677 6928
rect 9699 7013 9726 7021
rect 9699 6996 9704 7013
rect 9721 6996 9726 7013
rect 9699 6979 9726 6996
rect 9699 6962 9704 6979
rect 9721 6962 9726 6979
rect 9699 6945 9726 6962
rect 9699 6928 9704 6945
rect 9721 6928 9726 6945
rect 9699 6920 9726 6928
rect 10062 7013 10089 7021
rect 10062 6996 10067 7013
rect 10084 6996 10089 7013
rect 10062 6979 10089 6996
rect 10062 6962 10067 6979
rect 10084 6962 10089 6979
rect 10062 6945 10089 6962
rect 10062 6928 10067 6945
rect 10084 6928 10089 6945
rect 10062 6920 10089 6928
rect 10111 7013 10169 7021
rect 10111 6996 10147 7013
rect 10164 6996 10169 7013
rect 10111 6979 10169 6996
rect 10111 6962 10147 6979
rect 10164 6962 10169 6979
rect 10111 6945 10169 6962
rect 10111 6928 10147 6945
rect 10164 6928 10169 6945
rect 10111 6920 10169 6928
rect 10186 7013 10213 7021
rect 10186 6996 10191 7013
rect 10208 6996 10213 7013
rect 10186 6979 10213 6996
rect 10186 6962 10191 6979
rect 10208 6962 10213 6979
rect 10186 6945 10213 6962
rect 10186 6928 10191 6945
rect 10208 6928 10213 6945
rect 9575 6886 9579 6905
rect 9598 6886 9602 6905
rect 10186 6905 10213 6928
rect 10230 7013 10288 7021
rect 10230 6996 10235 7013
rect 10252 6996 10288 7013
rect 10230 6979 10288 6996
rect 10230 6962 10235 6979
rect 10252 6962 10288 6979
rect 10230 6945 10288 6962
rect 10230 6928 10235 6945
rect 10252 6928 10288 6945
rect 10230 6920 10288 6928
rect 10310 7013 10337 7021
rect 10310 6996 10315 7013
rect 10332 6996 10337 7013
rect 10310 6979 10337 6996
rect 10310 6962 10315 6979
rect 10332 6962 10337 6979
rect 10310 6945 10337 6962
rect 10310 6928 10315 6945
rect 10332 6928 10337 6945
rect 10310 6920 10337 6928
rect 10673 7013 10700 7021
rect 10673 6996 10678 7013
rect 10695 6996 10700 7013
rect 10673 6979 10700 6996
rect 10673 6962 10678 6979
rect 10695 6962 10700 6979
rect 10673 6945 10700 6962
rect 10673 6928 10678 6945
rect 10695 6928 10700 6945
rect 10673 6920 10700 6928
rect 10722 7013 10780 7021
rect 10722 6996 10758 7013
rect 10775 6996 10780 7013
rect 10722 6979 10780 6996
rect 10722 6962 10758 6979
rect 10775 6962 10780 6979
rect 10722 6945 10780 6962
rect 10722 6928 10758 6945
rect 10775 6928 10780 6945
rect 10722 6920 10780 6928
rect 10797 7013 10824 7021
rect 10797 6996 10802 7013
rect 10819 6996 10824 7013
rect 10797 6979 10824 6996
rect 10797 6962 10802 6979
rect 10819 6962 10824 6979
rect 10797 6945 10824 6962
rect 10797 6928 10802 6945
rect 10819 6928 10824 6945
rect 10186 6886 10190 6905
rect 10209 6886 10213 6905
rect 10797 6905 10824 6928
rect 10841 7013 10899 7021
rect 10841 6996 10846 7013
rect 10863 6996 10899 7013
rect 10841 6979 10899 6996
rect 10841 6962 10846 6979
rect 10863 6962 10899 6979
rect 10841 6945 10899 6962
rect 10841 6928 10846 6945
rect 10863 6928 10899 6945
rect 10841 6920 10899 6928
rect 10921 7013 10948 7021
rect 10921 6996 10926 7013
rect 10943 6996 10948 7013
rect 10921 6979 10948 6996
rect 10921 6962 10926 6979
rect 10943 6962 10948 6979
rect 10921 6945 10948 6962
rect 10921 6928 10926 6945
rect 10943 6928 10948 6945
rect 10921 6920 10948 6928
rect 11251 7013 11278 7021
rect 11251 6996 11256 7013
rect 11273 6996 11278 7013
rect 11251 6979 11278 6996
rect 11251 6962 11256 6979
rect 11273 6962 11278 6979
rect 11251 6945 11278 6962
rect 11251 6928 11256 6945
rect 11273 6928 11278 6945
rect 11251 6920 11278 6928
rect 11300 7013 11358 7021
rect 11300 6996 11336 7013
rect 11353 6996 11358 7013
rect 11300 6979 11358 6996
rect 11300 6962 11336 6979
rect 11353 6962 11358 6979
rect 11300 6945 11358 6962
rect 11300 6928 11336 6945
rect 11353 6928 11358 6945
rect 11300 6920 11358 6928
rect 11375 7013 11402 7021
rect 11375 6996 11380 7013
rect 11397 6996 11402 7013
rect 11375 6979 11402 6996
rect 11375 6962 11380 6979
rect 11397 6962 11402 6979
rect 11375 6945 11402 6962
rect 11375 6928 11380 6945
rect 11397 6928 11402 6945
rect 10797 6886 10801 6905
rect 10820 6886 10824 6905
rect 11375 6905 11402 6928
rect 11419 7013 11477 7021
rect 11419 6996 11424 7013
rect 11441 6996 11477 7013
rect 11419 6979 11477 6996
rect 11419 6962 11424 6979
rect 11441 6962 11477 6979
rect 11419 6945 11477 6962
rect 11419 6928 11424 6945
rect 11441 6928 11477 6945
rect 11419 6920 11477 6928
rect 11499 7013 11526 7021
rect 11499 6996 11504 7013
rect 11521 6996 11526 7013
rect 11499 6979 11526 6996
rect 11499 6962 11504 6979
rect 11521 6962 11526 6979
rect 11499 6945 11526 6962
rect 11499 6928 11504 6945
rect 11521 6928 11526 6945
rect 11499 6920 11526 6928
rect 11862 7013 11889 7021
rect 11862 6996 11867 7013
rect 11884 6996 11889 7013
rect 11862 6979 11889 6996
rect 11862 6962 11867 6979
rect 11884 6962 11889 6979
rect 11862 6945 11889 6962
rect 11862 6928 11867 6945
rect 11884 6928 11889 6945
rect 11862 6920 11889 6928
rect 11911 7013 11969 7021
rect 11911 6996 11947 7013
rect 11964 6996 11969 7013
rect 11911 6979 11969 6996
rect 11911 6962 11947 6979
rect 11964 6962 11969 6979
rect 11911 6945 11969 6962
rect 11911 6928 11947 6945
rect 11964 6928 11969 6945
rect 11911 6920 11969 6928
rect 11986 7013 12013 7021
rect 11986 6996 11991 7013
rect 12008 6996 12013 7013
rect 11986 6979 12013 6996
rect 11986 6962 11991 6979
rect 12008 6962 12013 6979
rect 11986 6945 12013 6962
rect 11986 6928 11991 6945
rect 12008 6928 12013 6945
rect 11375 6886 11379 6905
rect 11398 6886 11402 6905
rect 11986 6905 12013 6928
rect 12030 7013 12088 7021
rect 12030 6996 12035 7013
rect 12052 6996 12088 7013
rect 12030 6979 12088 6996
rect 12030 6962 12035 6979
rect 12052 6962 12088 6979
rect 12030 6945 12088 6962
rect 12030 6928 12035 6945
rect 12052 6928 12088 6945
rect 12030 6920 12088 6928
rect 12110 7013 12137 7021
rect 12110 6996 12115 7013
rect 12132 6996 12137 7013
rect 12110 6979 12137 6996
rect 12110 6962 12115 6979
rect 12132 6962 12137 6979
rect 12110 6945 12137 6962
rect 12110 6928 12115 6945
rect 12132 6928 12137 6945
rect 12110 6920 12137 6928
rect 12473 7013 12500 7021
rect 12473 6996 12478 7013
rect 12495 6996 12500 7013
rect 12473 6979 12500 6996
rect 12473 6962 12478 6979
rect 12495 6962 12500 6979
rect 12473 6945 12500 6962
rect 12473 6928 12478 6945
rect 12495 6928 12500 6945
rect 12473 6920 12500 6928
rect 12522 7013 12580 7021
rect 12522 6996 12558 7013
rect 12575 6996 12580 7013
rect 12522 6979 12580 6996
rect 12522 6962 12558 6979
rect 12575 6962 12580 6979
rect 12522 6945 12580 6962
rect 12522 6928 12558 6945
rect 12575 6928 12580 6945
rect 12522 6920 12580 6928
rect 12597 7013 12624 7021
rect 12597 6996 12602 7013
rect 12619 6996 12624 7013
rect 12597 6979 12624 6996
rect 12597 6962 12602 6979
rect 12619 6962 12624 6979
rect 12597 6945 12624 6962
rect 12597 6928 12602 6945
rect 12619 6928 12624 6945
rect 11986 6886 11990 6905
rect 12009 6886 12013 6905
rect 12597 6905 12624 6928
rect 12641 7013 12699 7021
rect 12641 6996 12646 7013
rect 12663 6996 12699 7013
rect 12641 6979 12699 6996
rect 12641 6962 12646 6979
rect 12663 6962 12699 6979
rect 12641 6945 12699 6962
rect 12641 6928 12646 6945
rect 12663 6928 12699 6945
rect 12641 6920 12699 6928
rect 12721 7013 12748 7021
rect 12721 6996 12726 7013
rect 12743 6996 12748 7013
rect 12721 6979 12748 6996
rect 12721 6962 12726 6979
rect 12743 6962 12748 6979
rect 12721 6945 12748 6962
rect 12721 6928 12726 6945
rect 12743 6928 12748 6945
rect 12721 6920 12748 6928
rect 12597 6886 12601 6905
rect 12620 6886 12624 6905
rect 9575 6772 9579 6791
rect 9598 6772 9602 6791
rect 9500 6749 9558 6757
rect 9500 6732 9536 6749
rect 9553 6732 9558 6749
rect 9500 6715 9558 6732
rect 9500 6698 9536 6715
rect 9553 6698 9558 6715
rect 9500 6681 9558 6698
rect 9500 6664 9536 6681
rect 9553 6664 9558 6681
rect 9500 6647 9558 6664
rect 9500 6630 9536 6647
rect 9553 6630 9558 6647
rect 9500 6613 9558 6630
rect 9500 6596 9536 6613
rect 9553 6596 9558 6613
rect 9500 6579 9558 6596
rect 9500 6562 9536 6579
rect 9553 6562 9558 6579
rect 9500 6554 9558 6562
rect 9575 6749 9602 6772
rect 10186 6772 10190 6791
rect 10209 6772 10213 6791
rect 9575 6732 9580 6749
rect 9597 6732 9602 6749
rect 9575 6715 9602 6732
rect 9575 6698 9580 6715
rect 9597 6698 9602 6715
rect 9575 6681 9602 6698
rect 9575 6664 9580 6681
rect 9597 6664 9602 6681
rect 9575 6647 9602 6664
rect 9575 6630 9580 6647
rect 9597 6630 9602 6647
rect 9575 6613 9602 6630
rect 9575 6596 9580 6613
rect 9597 6596 9602 6613
rect 9575 6579 9602 6596
rect 9575 6562 9580 6579
rect 9597 6562 9602 6579
rect 9575 6554 9602 6562
rect 9619 6749 9677 6757
rect 9619 6732 9624 6749
rect 9641 6732 9677 6749
rect 9619 6715 9677 6732
rect 9619 6698 9624 6715
rect 9641 6698 9677 6715
rect 9619 6681 9677 6698
rect 9619 6664 9624 6681
rect 9641 6664 9677 6681
rect 9619 6647 9677 6664
rect 9619 6630 9624 6647
rect 9641 6630 9677 6647
rect 9619 6613 9677 6630
rect 9619 6596 9624 6613
rect 9641 6596 9677 6613
rect 9619 6579 9677 6596
rect 9619 6562 9624 6579
rect 9641 6562 9677 6579
rect 9619 6554 9677 6562
rect 9450 6477 9483 6485
rect 9450 6460 9458 6477
rect 9475 6460 9483 6477
rect 9450 6452 9483 6460
rect 9500 6467 9527 6554
rect 9549 6529 9582 6537
rect 9549 6512 9557 6529
rect 9574 6521 9582 6529
rect 9650 6521 9677 6554
rect 9574 6512 9677 6521
rect 9549 6504 9677 6512
rect 9595 6475 9628 6483
rect 9595 6467 9603 6475
rect 9500 6458 9603 6467
rect 9620 6458 9628 6475
rect 9500 6450 9628 6458
rect 9450 6423 9483 6431
rect 9450 6406 9458 6423
rect 9475 6406 9483 6423
rect 9450 6398 9483 6406
rect 9500 6381 9527 6450
rect 9650 6381 9677 6504
rect 10111 6749 10169 6757
rect 10111 6732 10147 6749
rect 10164 6732 10169 6749
rect 10111 6715 10169 6732
rect 10111 6698 10147 6715
rect 10164 6698 10169 6715
rect 10111 6681 10169 6698
rect 10111 6664 10147 6681
rect 10164 6664 10169 6681
rect 10111 6647 10169 6664
rect 10111 6630 10147 6647
rect 10164 6630 10169 6647
rect 10111 6613 10169 6630
rect 10111 6596 10147 6613
rect 10164 6596 10169 6613
rect 10111 6579 10169 6596
rect 10111 6562 10147 6579
rect 10164 6562 10169 6579
rect 10111 6554 10169 6562
rect 10186 6749 10213 6772
rect 10797 6772 10801 6791
rect 10820 6772 10824 6791
rect 10186 6732 10191 6749
rect 10208 6732 10213 6749
rect 10186 6715 10213 6732
rect 10186 6698 10191 6715
rect 10208 6698 10213 6715
rect 10186 6681 10213 6698
rect 10186 6664 10191 6681
rect 10208 6664 10213 6681
rect 10186 6647 10213 6664
rect 10186 6630 10191 6647
rect 10208 6630 10213 6647
rect 10186 6613 10213 6630
rect 10186 6596 10191 6613
rect 10208 6596 10213 6613
rect 10186 6579 10213 6596
rect 10186 6562 10191 6579
rect 10208 6562 10213 6579
rect 10186 6554 10213 6562
rect 10230 6749 10288 6757
rect 10230 6732 10235 6749
rect 10252 6732 10288 6749
rect 10230 6715 10288 6732
rect 10230 6698 10235 6715
rect 10252 6698 10288 6715
rect 10230 6681 10288 6698
rect 10230 6664 10235 6681
rect 10252 6664 10288 6681
rect 10230 6647 10288 6664
rect 10230 6630 10235 6647
rect 10252 6630 10288 6647
rect 10230 6613 10288 6630
rect 10230 6596 10235 6613
rect 10252 6596 10288 6613
rect 10230 6579 10288 6596
rect 10230 6562 10235 6579
rect 10252 6562 10288 6579
rect 10230 6554 10288 6562
rect 10061 6477 10094 6485
rect 10061 6460 10069 6477
rect 10086 6460 10094 6477
rect 10061 6452 10094 6460
rect 10111 6467 10138 6554
rect 10160 6529 10193 6537
rect 10160 6512 10168 6529
rect 10185 6521 10193 6529
rect 10261 6521 10288 6554
rect 10185 6512 10288 6521
rect 10160 6504 10288 6512
rect 10206 6475 10239 6483
rect 10206 6467 10214 6475
rect 10111 6458 10214 6467
rect 10231 6458 10239 6475
rect 10111 6450 10239 6458
rect 9694 6439 9727 6447
rect 9694 6422 9702 6439
rect 9719 6422 9727 6439
rect 9694 6414 9727 6422
rect 10061 6423 10094 6431
rect 10061 6406 10069 6423
rect 10086 6406 10094 6423
rect 10061 6398 10094 6406
rect 10111 6381 10138 6450
rect 10261 6381 10288 6504
rect 10722 6749 10780 6757
rect 10722 6732 10758 6749
rect 10775 6732 10780 6749
rect 10722 6715 10780 6732
rect 10722 6698 10758 6715
rect 10775 6698 10780 6715
rect 10722 6681 10780 6698
rect 10722 6664 10758 6681
rect 10775 6664 10780 6681
rect 10722 6647 10780 6664
rect 10722 6630 10758 6647
rect 10775 6630 10780 6647
rect 10722 6613 10780 6630
rect 10722 6596 10758 6613
rect 10775 6596 10780 6613
rect 10722 6579 10780 6596
rect 10722 6562 10758 6579
rect 10775 6562 10780 6579
rect 10722 6554 10780 6562
rect 10797 6749 10824 6772
rect 11375 6772 11379 6791
rect 11398 6772 11402 6791
rect 10797 6732 10802 6749
rect 10819 6732 10824 6749
rect 10797 6715 10824 6732
rect 10797 6698 10802 6715
rect 10819 6698 10824 6715
rect 10797 6681 10824 6698
rect 10797 6664 10802 6681
rect 10819 6664 10824 6681
rect 10797 6647 10824 6664
rect 10797 6630 10802 6647
rect 10819 6630 10824 6647
rect 10797 6613 10824 6630
rect 10797 6596 10802 6613
rect 10819 6596 10824 6613
rect 10797 6579 10824 6596
rect 10797 6562 10802 6579
rect 10819 6562 10824 6579
rect 10797 6554 10824 6562
rect 10841 6749 10899 6757
rect 10841 6732 10846 6749
rect 10863 6732 10899 6749
rect 10841 6715 10899 6732
rect 10841 6698 10846 6715
rect 10863 6698 10899 6715
rect 10841 6681 10899 6698
rect 10841 6664 10846 6681
rect 10863 6664 10899 6681
rect 10841 6647 10899 6664
rect 10841 6630 10846 6647
rect 10863 6630 10899 6647
rect 10841 6613 10899 6630
rect 10841 6596 10846 6613
rect 10863 6596 10899 6613
rect 10841 6579 10899 6596
rect 10841 6562 10846 6579
rect 10863 6562 10899 6579
rect 10841 6554 10899 6562
rect 10672 6477 10705 6485
rect 10672 6460 10680 6477
rect 10697 6460 10705 6477
rect 10672 6452 10705 6460
rect 10722 6467 10749 6554
rect 10771 6529 10804 6537
rect 10771 6512 10779 6529
rect 10796 6521 10804 6529
rect 10872 6521 10899 6554
rect 10796 6512 10899 6521
rect 10771 6504 10899 6512
rect 10817 6475 10850 6483
rect 10817 6467 10825 6475
rect 10722 6458 10825 6467
rect 10842 6458 10850 6475
rect 10722 6450 10850 6458
rect 10305 6439 10338 6447
rect 10305 6422 10313 6439
rect 10330 6422 10338 6439
rect 10305 6414 10338 6422
rect 10672 6423 10705 6431
rect 10672 6406 10680 6423
rect 10697 6406 10705 6423
rect 10672 6398 10705 6406
rect 10722 6381 10749 6450
rect 10872 6381 10899 6504
rect 11300 6749 11358 6757
rect 11300 6732 11336 6749
rect 11353 6732 11358 6749
rect 11300 6715 11358 6732
rect 11300 6698 11336 6715
rect 11353 6698 11358 6715
rect 11300 6681 11358 6698
rect 11300 6664 11336 6681
rect 11353 6664 11358 6681
rect 11300 6647 11358 6664
rect 11300 6630 11336 6647
rect 11353 6630 11358 6647
rect 11300 6613 11358 6630
rect 11300 6596 11336 6613
rect 11353 6596 11358 6613
rect 11300 6579 11358 6596
rect 11300 6562 11336 6579
rect 11353 6562 11358 6579
rect 11300 6554 11358 6562
rect 11375 6749 11402 6772
rect 11986 6772 11990 6791
rect 12009 6772 12013 6791
rect 11375 6732 11380 6749
rect 11397 6732 11402 6749
rect 11375 6715 11402 6732
rect 11375 6698 11380 6715
rect 11397 6698 11402 6715
rect 11375 6681 11402 6698
rect 11375 6664 11380 6681
rect 11397 6664 11402 6681
rect 11375 6647 11402 6664
rect 11375 6630 11380 6647
rect 11397 6630 11402 6647
rect 11375 6613 11402 6630
rect 11375 6596 11380 6613
rect 11397 6596 11402 6613
rect 11375 6579 11402 6596
rect 11375 6562 11380 6579
rect 11397 6562 11402 6579
rect 11375 6554 11402 6562
rect 11419 6749 11477 6757
rect 11419 6732 11424 6749
rect 11441 6732 11477 6749
rect 11419 6715 11477 6732
rect 11419 6698 11424 6715
rect 11441 6698 11477 6715
rect 11419 6681 11477 6698
rect 11419 6664 11424 6681
rect 11441 6664 11477 6681
rect 11419 6647 11477 6664
rect 11419 6630 11424 6647
rect 11441 6630 11477 6647
rect 11419 6613 11477 6630
rect 11419 6596 11424 6613
rect 11441 6596 11477 6613
rect 11419 6579 11477 6596
rect 11419 6562 11424 6579
rect 11441 6562 11477 6579
rect 11419 6554 11477 6562
rect 11250 6477 11283 6485
rect 11250 6460 11258 6477
rect 11275 6460 11283 6477
rect 11250 6452 11283 6460
rect 11300 6467 11327 6554
rect 11349 6529 11382 6537
rect 11349 6512 11357 6529
rect 11374 6521 11382 6529
rect 11450 6521 11477 6554
rect 11374 6512 11477 6521
rect 11349 6504 11477 6512
rect 11395 6475 11428 6483
rect 11395 6467 11403 6475
rect 11300 6458 11403 6467
rect 11420 6458 11428 6475
rect 11300 6450 11428 6458
rect 10916 6439 10949 6447
rect 10916 6422 10924 6439
rect 10941 6422 10949 6439
rect 10916 6414 10949 6422
rect 11250 6423 11283 6431
rect 11250 6406 11258 6423
rect 11275 6406 11283 6423
rect 11250 6398 11283 6406
rect 11300 6381 11327 6450
rect 11450 6381 11477 6504
rect 11911 6749 11969 6757
rect 11911 6732 11947 6749
rect 11964 6732 11969 6749
rect 11911 6715 11969 6732
rect 11911 6698 11947 6715
rect 11964 6698 11969 6715
rect 11911 6681 11969 6698
rect 11911 6664 11947 6681
rect 11964 6664 11969 6681
rect 11911 6647 11969 6664
rect 11911 6630 11947 6647
rect 11964 6630 11969 6647
rect 11911 6613 11969 6630
rect 11911 6596 11947 6613
rect 11964 6596 11969 6613
rect 11911 6579 11969 6596
rect 11911 6562 11947 6579
rect 11964 6562 11969 6579
rect 11911 6554 11969 6562
rect 11986 6749 12013 6772
rect 12597 6772 12601 6791
rect 12620 6772 12624 6791
rect 11986 6732 11991 6749
rect 12008 6732 12013 6749
rect 11986 6715 12013 6732
rect 11986 6698 11991 6715
rect 12008 6698 12013 6715
rect 11986 6681 12013 6698
rect 11986 6664 11991 6681
rect 12008 6664 12013 6681
rect 11986 6647 12013 6664
rect 11986 6630 11991 6647
rect 12008 6630 12013 6647
rect 11986 6613 12013 6630
rect 11986 6596 11991 6613
rect 12008 6596 12013 6613
rect 11986 6579 12013 6596
rect 11986 6562 11991 6579
rect 12008 6562 12013 6579
rect 11986 6554 12013 6562
rect 12030 6749 12088 6757
rect 12030 6732 12035 6749
rect 12052 6732 12088 6749
rect 12030 6715 12088 6732
rect 12030 6698 12035 6715
rect 12052 6698 12088 6715
rect 12030 6681 12088 6698
rect 12030 6664 12035 6681
rect 12052 6664 12088 6681
rect 12030 6647 12088 6664
rect 12030 6630 12035 6647
rect 12052 6630 12088 6647
rect 12030 6613 12088 6630
rect 12030 6596 12035 6613
rect 12052 6596 12088 6613
rect 12030 6579 12088 6596
rect 12030 6562 12035 6579
rect 12052 6562 12088 6579
rect 12030 6554 12088 6562
rect 11861 6477 11894 6485
rect 11861 6460 11869 6477
rect 11886 6460 11894 6477
rect 11861 6452 11894 6460
rect 11911 6467 11938 6554
rect 11960 6529 11993 6537
rect 11960 6512 11968 6529
rect 11985 6521 11993 6529
rect 12061 6521 12088 6554
rect 11985 6512 12088 6521
rect 11960 6504 12088 6512
rect 12006 6475 12039 6483
rect 12006 6467 12014 6475
rect 11911 6458 12014 6467
rect 12031 6458 12039 6475
rect 11911 6450 12039 6458
rect 11494 6439 11527 6447
rect 11494 6422 11502 6439
rect 11519 6422 11527 6439
rect 11494 6414 11527 6422
rect 11861 6423 11894 6431
rect 11861 6406 11869 6423
rect 11886 6406 11894 6423
rect 11861 6398 11894 6406
rect 11911 6381 11938 6450
rect 12061 6381 12088 6504
rect 12522 6749 12580 6757
rect 12522 6732 12558 6749
rect 12575 6732 12580 6749
rect 12522 6715 12580 6732
rect 12522 6698 12558 6715
rect 12575 6698 12580 6715
rect 12522 6681 12580 6698
rect 12522 6664 12558 6681
rect 12575 6664 12580 6681
rect 12522 6647 12580 6664
rect 12522 6630 12558 6647
rect 12575 6630 12580 6647
rect 12522 6613 12580 6630
rect 12522 6596 12558 6613
rect 12575 6596 12580 6613
rect 12522 6579 12580 6596
rect 12522 6562 12558 6579
rect 12575 6562 12580 6579
rect 12522 6554 12580 6562
rect 12597 6749 12624 6772
rect 12597 6732 12602 6749
rect 12619 6732 12624 6749
rect 12597 6715 12624 6732
rect 12597 6698 12602 6715
rect 12619 6698 12624 6715
rect 12597 6681 12624 6698
rect 12597 6664 12602 6681
rect 12619 6664 12624 6681
rect 12597 6647 12624 6664
rect 12597 6630 12602 6647
rect 12619 6630 12624 6647
rect 12597 6613 12624 6630
rect 12597 6596 12602 6613
rect 12619 6596 12624 6613
rect 12597 6579 12624 6596
rect 12597 6562 12602 6579
rect 12619 6562 12624 6579
rect 12597 6554 12624 6562
rect 12641 6749 12699 6757
rect 12641 6732 12646 6749
rect 12663 6732 12699 6749
rect 12641 6715 12699 6732
rect 12641 6698 12646 6715
rect 12663 6698 12699 6715
rect 12641 6681 12699 6698
rect 12641 6664 12646 6681
rect 12663 6664 12699 6681
rect 12641 6647 12699 6664
rect 12641 6630 12646 6647
rect 12663 6630 12699 6647
rect 12641 6613 12699 6630
rect 12641 6596 12646 6613
rect 12663 6596 12699 6613
rect 12641 6579 12699 6596
rect 12641 6562 12646 6579
rect 12663 6562 12699 6579
rect 12641 6554 12699 6562
rect 12472 6477 12505 6485
rect 12472 6460 12480 6477
rect 12497 6460 12505 6477
rect 12472 6452 12505 6460
rect 12522 6467 12549 6554
rect 12571 6529 12604 6537
rect 12571 6512 12579 6529
rect 12596 6521 12604 6529
rect 12672 6521 12699 6554
rect 12596 6512 12699 6521
rect 12571 6504 12699 6512
rect 12617 6475 12650 6483
rect 12617 6467 12625 6475
rect 12522 6458 12625 6467
rect 12642 6458 12650 6475
rect 12522 6450 12650 6458
rect 12105 6439 12138 6447
rect 12105 6422 12113 6439
rect 12130 6422 12138 6439
rect 12105 6414 12138 6422
rect 12472 6423 12505 6431
rect 12472 6406 12480 6423
rect 12497 6406 12505 6423
rect 12472 6398 12505 6406
rect 12522 6381 12549 6450
rect 12672 6381 12699 6504
rect 12716 6439 12749 6447
rect 12716 6422 12724 6439
rect 12741 6422 12749 6439
rect 12716 6414 12749 6422
rect 9451 6373 9478 6381
rect 9451 6356 9456 6373
rect 9473 6356 9478 6373
rect 9451 6339 9478 6356
rect 9451 6322 9456 6339
rect 9473 6322 9478 6339
rect 9451 6305 9478 6322
rect 9451 6288 9456 6305
rect 9473 6288 9478 6305
rect 9451 6280 9478 6288
rect 9500 6373 9558 6381
rect 9500 6356 9536 6373
rect 9553 6356 9558 6373
rect 9500 6339 9558 6356
rect 9500 6322 9536 6339
rect 9553 6322 9558 6339
rect 9500 6305 9558 6322
rect 9500 6288 9536 6305
rect 9553 6288 9558 6305
rect 9500 6280 9558 6288
rect 9575 6373 9602 6381
rect 9575 6356 9580 6373
rect 9597 6356 9602 6373
rect 9575 6339 9602 6356
rect 9575 6322 9580 6339
rect 9597 6322 9602 6339
rect 9575 6305 9602 6322
rect 9575 6288 9580 6305
rect 9597 6288 9602 6305
rect 9575 6265 9602 6288
rect 9619 6373 9677 6381
rect 9619 6356 9624 6373
rect 9641 6356 9677 6373
rect 9619 6339 9677 6356
rect 9619 6322 9624 6339
rect 9641 6322 9677 6339
rect 9619 6305 9677 6322
rect 9619 6288 9624 6305
rect 9641 6288 9677 6305
rect 9619 6280 9677 6288
rect 9699 6373 9726 6381
rect 9699 6356 9704 6373
rect 9721 6356 9726 6373
rect 9699 6339 9726 6356
rect 9699 6322 9704 6339
rect 9721 6322 9726 6339
rect 9699 6305 9726 6322
rect 9699 6288 9704 6305
rect 9721 6288 9726 6305
rect 9699 6280 9726 6288
rect 10062 6373 10089 6381
rect 10062 6356 10067 6373
rect 10084 6356 10089 6373
rect 10062 6339 10089 6356
rect 10062 6322 10067 6339
rect 10084 6322 10089 6339
rect 10062 6305 10089 6322
rect 10062 6288 10067 6305
rect 10084 6288 10089 6305
rect 10062 6280 10089 6288
rect 10111 6373 10169 6381
rect 10111 6356 10147 6373
rect 10164 6356 10169 6373
rect 10111 6339 10169 6356
rect 10111 6322 10147 6339
rect 10164 6322 10169 6339
rect 10111 6305 10169 6322
rect 10111 6288 10147 6305
rect 10164 6288 10169 6305
rect 10111 6280 10169 6288
rect 10186 6373 10213 6381
rect 10186 6356 10191 6373
rect 10208 6356 10213 6373
rect 10186 6339 10213 6356
rect 10186 6322 10191 6339
rect 10208 6322 10213 6339
rect 10186 6305 10213 6322
rect 10186 6288 10191 6305
rect 10208 6288 10213 6305
rect 9575 6246 9579 6265
rect 9598 6246 9602 6265
rect 10186 6265 10213 6288
rect 10230 6373 10288 6381
rect 10230 6356 10235 6373
rect 10252 6356 10288 6373
rect 10230 6339 10288 6356
rect 10230 6322 10235 6339
rect 10252 6322 10288 6339
rect 10230 6305 10288 6322
rect 10230 6288 10235 6305
rect 10252 6288 10288 6305
rect 10230 6280 10288 6288
rect 10310 6373 10337 6381
rect 10310 6356 10315 6373
rect 10332 6356 10337 6373
rect 10310 6339 10337 6356
rect 10310 6322 10315 6339
rect 10332 6322 10337 6339
rect 10310 6305 10337 6322
rect 10310 6288 10315 6305
rect 10332 6288 10337 6305
rect 10310 6280 10337 6288
rect 10673 6373 10700 6381
rect 10673 6356 10678 6373
rect 10695 6356 10700 6373
rect 10673 6339 10700 6356
rect 10673 6322 10678 6339
rect 10695 6322 10700 6339
rect 10673 6305 10700 6322
rect 10673 6288 10678 6305
rect 10695 6288 10700 6305
rect 10673 6280 10700 6288
rect 10722 6373 10780 6381
rect 10722 6356 10758 6373
rect 10775 6356 10780 6373
rect 10722 6339 10780 6356
rect 10722 6322 10758 6339
rect 10775 6322 10780 6339
rect 10722 6305 10780 6322
rect 10722 6288 10758 6305
rect 10775 6288 10780 6305
rect 10722 6280 10780 6288
rect 10797 6373 10824 6381
rect 10797 6356 10802 6373
rect 10819 6356 10824 6373
rect 10797 6339 10824 6356
rect 10797 6322 10802 6339
rect 10819 6322 10824 6339
rect 10797 6305 10824 6322
rect 10797 6288 10802 6305
rect 10819 6288 10824 6305
rect 10186 6246 10190 6265
rect 10209 6246 10213 6265
rect 10797 6265 10824 6288
rect 10841 6373 10899 6381
rect 10841 6356 10846 6373
rect 10863 6356 10899 6373
rect 10841 6339 10899 6356
rect 10841 6322 10846 6339
rect 10863 6322 10899 6339
rect 10841 6305 10899 6322
rect 10841 6288 10846 6305
rect 10863 6288 10899 6305
rect 10841 6280 10899 6288
rect 10921 6373 10948 6381
rect 10921 6356 10926 6373
rect 10943 6356 10948 6373
rect 10921 6339 10948 6356
rect 10921 6322 10926 6339
rect 10943 6322 10948 6339
rect 10921 6305 10948 6322
rect 10921 6288 10926 6305
rect 10943 6288 10948 6305
rect 10921 6280 10948 6288
rect 11251 6373 11278 6381
rect 11251 6356 11256 6373
rect 11273 6356 11278 6373
rect 11251 6339 11278 6356
rect 11251 6322 11256 6339
rect 11273 6322 11278 6339
rect 11251 6305 11278 6322
rect 11251 6288 11256 6305
rect 11273 6288 11278 6305
rect 11251 6280 11278 6288
rect 11300 6373 11358 6381
rect 11300 6356 11336 6373
rect 11353 6356 11358 6373
rect 11300 6339 11358 6356
rect 11300 6322 11336 6339
rect 11353 6322 11358 6339
rect 11300 6305 11358 6322
rect 11300 6288 11336 6305
rect 11353 6288 11358 6305
rect 11300 6280 11358 6288
rect 11375 6373 11402 6381
rect 11375 6356 11380 6373
rect 11397 6356 11402 6373
rect 11375 6339 11402 6356
rect 11375 6322 11380 6339
rect 11397 6322 11402 6339
rect 11375 6305 11402 6322
rect 11375 6288 11380 6305
rect 11397 6288 11402 6305
rect 10797 6246 10801 6265
rect 10820 6246 10824 6265
rect 11375 6265 11402 6288
rect 11419 6373 11477 6381
rect 11419 6356 11424 6373
rect 11441 6356 11477 6373
rect 11419 6339 11477 6356
rect 11419 6322 11424 6339
rect 11441 6322 11477 6339
rect 11419 6305 11477 6322
rect 11419 6288 11424 6305
rect 11441 6288 11477 6305
rect 11419 6280 11477 6288
rect 11499 6373 11526 6381
rect 11499 6356 11504 6373
rect 11521 6356 11526 6373
rect 11499 6339 11526 6356
rect 11499 6322 11504 6339
rect 11521 6322 11526 6339
rect 11499 6305 11526 6322
rect 11499 6288 11504 6305
rect 11521 6288 11526 6305
rect 11499 6280 11526 6288
rect 11862 6373 11889 6381
rect 11862 6356 11867 6373
rect 11884 6356 11889 6373
rect 11862 6339 11889 6356
rect 11862 6322 11867 6339
rect 11884 6322 11889 6339
rect 11862 6305 11889 6322
rect 11862 6288 11867 6305
rect 11884 6288 11889 6305
rect 11862 6280 11889 6288
rect 11911 6373 11969 6381
rect 11911 6356 11947 6373
rect 11964 6356 11969 6373
rect 11911 6339 11969 6356
rect 11911 6322 11947 6339
rect 11964 6322 11969 6339
rect 11911 6305 11969 6322
rect 11911 6288 11947 6305
rect 11964 6288 11969 6305
rect 11911 6280 11969 6288
rect 11986 6373 12013 6381
rect 11986 6356 11991 6373
rect 12008 6356 12013 6373
rect 11986 6339 12013 6356
rect 11986 6322 11991 6339
rect 12008 6322 12013 6339
rect 11986 6305 12013 6322
rect 11986 6288 11991 6305
rect 12008 6288 12013 6305
rect 11375 6246 11379 6265
rect 11398 6246 11402 6265
rect 11986 6265 12013 6288
rect 12030 6373 12088 6381
rect 12030 6356 12035 6373
rect 12052 6356 12088 6373
rect 12030 6339 12088 6356
rect 12030 6322 12035 6339
rect 12052 6322 12088 6339
rect 12030 6305 12088 6322
rect 12030 6288 12035 6305
rect 12052 6288 12088 6305
rect 12030 6280 12088 6288
rect 12110 6373 12137 6381
rect 12110 6356 12115 6373
rect 12132 6356 12137 6373
rect 12110 6339 12137 6356
rect 12110 6322 12115 6339
rect 12132 6322 12137 6339
rect 12110 6305 12137 6322
rect 12110 6288 12115 6305
rect 12132 6288 12137 6305
rect 12110 6280 12137 6288
rect 12473 6373 12500 6381
rect 12473 6356 12478 6373
rect 12495 6356 12500 6373
rect 12473 6339 12500 6356
rect 12473 6322 12478 6339
rect 12495 6322 12500 6339
rect 12473 6305 12500 6322
rect 12473 6288 12478 6305
rect 12495 6288 12500 6305
rect 12473 6280 12500 6288
rect 12522 6373 12580 6381
rect 12522 6356 12558 6373
rect 12575 6356 12580 6373
rect 12522 6339 12580 6356
rect 12522 6322 12558 6339
rect 12575 6322 12580 6339
rect 12522 6305 12580 6322
rect 12522 6288 12558 6305
rect 12575 6288 12580 6305
rect 12522 6280 12580 6288
rect 12597 6373 12624 6381
rect 12597 6356 12602 6373
rect 12619 6356 12624 6373
rect 12597 6339 12624 6356
rect 12597 6322 12602 6339
rect 12619 6322 12624 6339
rect 12597 6305 12624 6322
rect 12597 6288 12602 6305
rect 12619 6288 12624 6305
rect 11986 6246 11990 6265
rect 12009 6246 12013 6265
rect 12597 6265 12624 6288
rect 12641 6373 12699 6381
rect 12641 6356 12646 6373
rect 12663 6356 12699 6373
rect 12641 6339 12699 6356
rect 12641 6322 12646 6339
rect 12663 6322 12699 6339
rect 12641 6305 12699 6322
rect 12641 6288 12646 6305
rect 12663 6288 12699 6305
rect 12641 6280 12699 6288
rect 12721 6373 12748 6381
rect 12721 6356 12726 6373
rect 12743 6356 12748 6373
rect 12721 6339 12748 6356
rect 12721 6322 12726 6339
rect 12743 6322 12748 6339
rect 12721 6305 12748 6322
rect 12721 6288 12726 6305
rect 12743 6288 12748 6305
rect 12721 6280 12748 6288
rect 12597 6246 12601 6265
rect 12620 6246 12624 6265
rect 9575 6122 9579 6141
rect 9598 6122 9602 6141
rect 9500 6099 9558 6107
rect 9500 6082 9536 6099
rect 9553 6082 9558 6099
rect 9500 6065 9558 6082
rect 9500 6048 9536 6065
rect 9553 6048 9558 6065
rect 9500 6031 9558 6048
rect 9500 6014 9536 6031
rect 9553 6014 9558 6031
rect 9500 5997 9558 6014
rect 9500 5980 9536 5997
rect 9553 5980 9558 5997
rect 9500 5963 9558 5980
rect 9500 5946 9536 5963
rect 9553 5946 9558 5963
rect 9500 5929 9558 5946
rect 9500 5912 9536 5929
rect 9553 5912 9558 5929
rect 9500 5904 9558 5912
rect 9575 6099 9602 6122
rect 10186 6122 10190 6141
rect 10209 6122 10213 6141
rect 9575 6082 9580 6099
rect 9597 6082 9602 6099
rect 9575 6065 9602 6082
rect 9575 6048 9580 6065
rect 9597 6048 9602 6065
rect 9575 6031 9602 6048
rect 9575 6014 9580 6031
rect 9597 6014 9602 6031
rect 9575 5997 9602 6014
rect 9575 5980 9580 5997
rect 9597 5980 9602 5997
rect 9575 5963 9602 5980
rect 9575 5946 9580 5963
rect 9597 5946 9602 5963
rect 9575 5929 9602 5946
rect 9575 5912 9580 5929
rect 9597 5912 9602 5929
rect 9575 5904 9602 5912
rect 9619 6099 9677 6107
rect 9619 6082 9624 6099
rect 9641 6082 9677 6099
rect 9619 6065 9677 6082
rect 9619 6048 9624 6065
rect 9641 6048 9677 6065
rect 9619 6031 9677 6048
rect 9619 6014 9624 6031
rect 9641 6014 9677 6031
rect 9619 5997 9677 6014
rect 9619 5980 9624 5997
rect 9641 5980 9677 5997
rect 9619 5963 9677 5980
rect 9619 5946 9624 5963
rect 9641 5946 9677 5963
rect 9619 5929 9677 5946
rect 9619 5912 9624 5929
rect 9641 5912 9677 5929
rect 9619 5904 9677 5912
rect 9450 5827 9483 5835
rect 9450 5810 9458 5827
rect 9475 5810 9483 5827
rect 9450 5802 9483 5810
rect 9500 5817 9527 5904
rect 9549 5879 9582 5887
rect 9549 5862 9557 5879
rect 9574 5871 9582 5879
rect 9650 5871 9677 5904
rect 9574 5862 9677 5871
rect 9549 5854 9677 5862
rect 9595 5825 9628 5833
rect 9595 5817 9603 5825
rect 9500 5808 9603 5817
rect 9620 5808 9628 5825
rect 9500 5800 9628 5808
rect 9450 5773 9483 5781
rect 9450 5756 9458 5773
rect 9475 5756 9483 5773
rect 9450 5748 9483 5756
rect 9500 5731 9527 5800
rect 9650 5731 9677 5854
rect 10111 6099 10169 6107
rect 10111 6082 10147 6099
rect 10164 6082 10169 6099
rect 10111 6065 10169 6082
rect 10111 6048 10147 6065
rect 10164 6048 10169 6065
rect 10111 6031 10169 6048
rect 10111 6014 10147 6031
rect 10164 6014 10169 6031
rect 10111 5997 10169 6014
rect 10111 5980 10147 5997
rect 10164 5980 10169 5997
rect 10111 5963 10169 5980
rect 10111 5946 10147 5963
rect 10164 5946 10169 5963
rect 10111 5929 10169 5946
rect 10111 5912 10147 5929
rect 10164 5912 10169 5929
rect 10111 5904 10169 5912
rect 10186 6099 10213 6122
rect 10797 6122 10801 6141
rect 10820 6122 10824 6141
rect 10186 6082 10191 6099
rect 10208 6082 10213 6099
rect 10186 6065 10213 6082
rect 10186 6048 10191 6065
rect 10208 6048 10213 6065
rect 10186 6031 10213 6048
rect 10186 6014 10191 6031
rect 10208 6014 10213 6031
rect 10186 5997 10213 6014
rect 10186 5980 10191 5997
rect 10208 5980 10213 5997
rect 10186 5963 10213 5980
rect 10186 5946 10191 5963
rect 10208 5946 10213 5963
rect 10186 5929 10213 5946
rect 10186 5912 10191 5929
rect 10208 5912 10213 5929
rect 10186 5904 10213 5912
rect 10230 6099 10288 6107
rect 10230 6082 10235 6099
rect 10252 6082 10288 6099
rect 10230 6065 10288 6082
rect 10230 6048 10235 6065
rect 10252 6048 10288 6065
rect 10230 6031 10288 6048
rect 10230 6014 10235 6031
rect 10252 6014 10288 6031
rect 10230 5997 10288 6014
rect 10230 5980 10235 5997
rect 10252 5980 10288 5997
rect 10230 5963 10288 5980
rect 10230 5946 10235 5963
rect 10252 5946 10288 5963
rect 10230 5929 10288 5946
rect 10230 5912 10235 5929
rect 10252 5912 10288 5929
rect 10230 5904 10288 5912
rect 10061 5827 10094 5835
rect 10061 5810 10069 5827
rect 10086 5810 10094 5827
rect 10061 5802 10094 5810
rect 10111 5817 10138 5904
rect 10160 5879 10193 5887
rect 10160 5862 10168 5879
rect 10185 5871 10193 5879
rect 10261 5871 10288 5904
rect 10185 5862 10288 5871
rect 10160 5854 10288 5862
rect 10206 5825 10239 5833
rect 10206 5817 10214 5825
rect 10111 5808 10214 5817
rect 10231 5808 10239 5825
rect 10111 5800 10239 5808
rect 9694 5789 9727 5797
rect 9694 5772 9702 5789
rect 9719 5772 9727 5789
rect 9694 5764 9727 5772
rect 10061 5773 10094 5781
rect 10061 5756 10069 5773
rect 10086 5756 10094 5773
rect 10061 5748 10094 5756
rect 10111 5731 10138 5800
rect 10261 5731 10288 5854
rect 10722 6099 10780 6107
rect 10722 6082 10758 6099
rect 10775 6082 10780 6099
rect 10722 6065 10780 6082
rect 10722 6048 10758 6065
rect 10775 6048 10780 6065
rect 10722 6031 10780 6048
rect 10722 6014 10758 6031
rect 10775 6014 10780 6031
rect 10722 5997 10780 6014
rect 10722 5980 10758 5997
rect 10775 5980 10780 5997
rect 10722 5963 10780 5980
rect 10722 5946 10758 5963
rect 10775 5946 10780 5963
rect 10722 5929 10780 5946
rect 10722 5912 10758 5929
rect 10775 5912 10780 5929
rect 10722 5904 10780 5912
rect 10797 6099 10824 6122
rect 11375 6122 11379 6141
rect 11398 6122 11402 6141
rect 10797 6082 10802 6099
rect 10819 6082 10824 6099
rect 10797 6065 10824 6082
rect 10797 6048 10802 6065
rect 10819 6048 10824 6065
rect 10797 6031 10824 6048
rect 10797 6014 10802 6031
rect 10819 6014 10824 6031
rect 10797 5997 10824 6014
rect 10797 5980 10802 5997
rect 10819 5980 10824 5997
rect 10797 5963 10824 5980
rect 10797 5946 10802 5963
rect 10819 5946 10824 5963
rect 10797 5929 10824 5946
rect 10797 5912 10802 5929
rect 10819 5912 10824 5929
rect 10797 5904 10824 5912
rect 10841 6099 10899 6107
rect 10841 6082 10846 6099
rect 10863 6082 10899 6099
rect 10841 6065 10899 6082
rect 10841 6048 10846 6065
rect 10863 6048 10899 6065
rect 10841 6031 10899 6048
rect 10841 6014 10846 6031
rect 10863 6014 10899 6031
rect 10841 5997 10899 6014
rect 10841 5980 10846 5997
rect 10863 5980 10899 5997
rect 10841 5963 10899 5980
rect 10841 5946 10846 5963
rect 10863 5946 10899 5963
rect 10841 5929 10899 5946
rect 10841 5912 10846 5929
rect 10863 5912 10899 5929
rect 10841 5904 10899 5912
rect 10672 5827 10705 5835
rect 10672 5810 10680 5827
rect 10697 5810 10705 5827
rect 10672 5802 10705 5810
rect 10722 5817 10749 5904
rect 10771 5879 10804 5887
rect 10771 5862 10779 5879
rect 10796 5871 10804 5879
rect 10872 5871 10899 5904
rect 10796 5862 10899 5871
rect 10771 5854 10899 5862
rect 10817 5825 10850 5833
rect 10817 5817 10825 5825
rect 10722 5808 10825 5817
rect 10842 5808 10850 5825
rect 10722 5800 10850 5808
rect 10305 5789 10338 5797
rect 10305 5772 10313 5789
rect 10330 5772 10338 5789
rect 10305 5764 10338 5772
rect 10672 5773 10705 5781
rect 10672 5756 10680 5773
rect 10697 5756 10705 5773
rect 10672 5748 10705 5756
rect 10722 5731 10749 5800
rect 10872 5731 10899 5854
rect 11300 6099 11358 6107
rect 11300 6082 11336 6099
rect 11353 6082 11358 6099
rect 11300 6065 11358 6082
rect 11300 6048 11336 6065
rect 11353 6048 11358 6065
rect 11300 6031 11358 6048
rect 11300 6014 11336 6031
rect 11353 6014 11358 6031
rect 11300 5997 11358 6014
rect 11300 5980 11336 5997
rect 11353 5980 11358 5997
rect 11300 5963 11358 5980
rect 11300 5946 11336 5963
rect 11353 5946 11358 5963
rect 11300 5929 11358 5946
rect 11300 5912 11336 5929
rect 11353 5912 11358 5929
rect 11300 5904 11358 5912
rect 11375 6099 11402 6122
rect 11986 6122 11990 6141
rect 12009 6122 12013 6141
rect 11375 6082 11380 6099
rect 11397 6082 11402 6099
rect 11375 6065 11402 6082
rect 11375 6048 11380 6065
rect 11397 6048 11402 6065
rect 11375 6031 11402 6048
rect 11375 6014 11380 6031
rect 11397 6014 11402 6031
rect 11375 5997 11402 6014
rect 11375 5980 11380 5997
rect 11397 5980 11402 5997
rect 11375 5963 11402 5980
rect 11375 5946 11380 5963
rect 11397 5946 11402 5963
rect 11375 5929 11402 5946
rect 11375 5912 11380 5929
rect 11397 5912 11402 5929
rect 11375 5904 11402 5912
rect 11419 6099 11477 6107
rect 11419 6082 11424 6099
rect 11441 6082 11477 6099
rect 11419 6065 11477 6082
rect 11419 6048 11424 6065
rect 11441 6048 11477 6065
rect 11419 6031 11477 6048
rect 11419 6014 11424 6031
rect 11441 6014 11477 6031
rect 11419 5997 11477 6014
rect 11419 5980 11424 5997
rect 11441 5980 11477 5997
rect 11419 5963 11477 5980
rect 11419 5946 11424 5963
rect 11441 5946 11477 5963
rect 11419 5929 11477 5946
rect 11419 5912 11424 5929
rect 11441 5912 11477 5929
rect 11419 5904 11477 5912
rect 11250 5827 11283 5835
rect 11250 5810 11258 5827
rect 11275 5810 11283 5827
rect 11250 5802 11283 5810
rect 11300 5817 11327 5904
rect 11349 5879 11382 5887
rect 11349 5862 11357 5879
rect 11374 5871 11382 5879
rect 11450 5871 11477 5904
rect 11374 5862 11477 5871
rect 11349 5854 11477 5862
rect 11395 5825 11428 5833
rect 11395 5817 11403 5825
rect 11300 5808 11403 5817
rect 11420 5808 11428 5825
rect 11300 5800 11428 5808
rect 10916 5789 10949 5797
rect 10916 5772 10924 5789
rect 10941 5772 10949 5789
rect 10916 5764 10949 5772
rect 11250 5773 11283 5781
rect 11250 5756 11258 5773
rect 11275 5756 11283 5773
rect 11250 5748 11283 5756
rect 11300 5731 11327 5800
rect 11450 5731 11477 5854
rect 11911 6099 11969 6107
rect 11911 6082 11947 6099
rect 11964 6082 11969 6099
rect 11911 6065 11969 6082
rect 11911 6048 11947 6065
rect 11964 6048 11969 6065
rect 11911 6031 11969 6048
rect 11911 6014 11947 6031
rect 11964 6014 11969 6031
rect 11911 5997 11969 6014
rect 11911 5980 11947 5997
rect 11964 5980 11969 5997
rect 11911 5963 11969 5980
rect 11911 5946 11947 5963
rect 11964 5946 11969 5963
rect 11911 5929 11969 5946
rect 11911 5912 11947 5929
rect 11964 5912 11969 5929
rect 11911 5904 11969 5912
rect 11986 6099 12013 6122
rect 12597 6122 12601 6141
rect 12620 6122 12624 6141
rect 11986 6082 11991 6099
rect 12008 6082 12013 6099
rect 11986 6065 12013 6082
rect 11986 6048 11991 6065
rect 12008 6048 12013 6065
rect 11986 6031 12013 6048
rect 11986 6014 11991 6031
rect 12008 6014 12013 6031
rect 11986 5997 12013 6014
rect 11986 5980 11991 5997
rect 12008 5980 12013 5997
rect 11986 5963 12013 5980
rect 11986 5946 11991 5963
rect 12008 5946 12013 5963
rect 11986 5929 12013 5946
rect 11986 5912 11991 5929
rect 12008 5912 12013 5929
rect 11986 5904 12013 5912
rect 12030 6099 12088 6107
rect 12030 6082 12035 6099
rect 12052 6082 12088 6099
rect 12030 6065 12088 6082
rect 12030 6048 12035 6065
rect 12052 6048 12088 6065
rect 12030 6031 12088 6048
rect 12030 6014 12035 6031
rect 12052 6014 12088 6031
rect 12030 5997 12088 6014
rect 12030 5980 12035 5997
rect 12052 5980 12088 5997
rect 12030 5963 12088 5980
rect 12030 5946 12035 5963
rect 12052 5946 12088 5963
rect 12030 5929 12088 5946
rect 12030 5912 12035 5929
rect 12052 5912 12088 5929
rect 12030 5904 12088 5912
rect 11861 5827 11894 5835
rect 11861 5810 11869 5827
rect 11886 5810 11894 5827
rect 11861 5802 11894 5810
rect 11911 5817 11938 5904
rect 11960 5879 11993 5887
rect 11960 5862 11968 5879
rect 11985 5871 11993 5879
rect 12061 5871 12088 5904
rect 11985 5862 12088 5871
rect 11960 5854 12088 5862
rect 12006 5825 12039 5833
rect 12006 5817 12014 5825
rect 11911 5808 12014 5817
rect 12031 5808 12039 5825
rect 11911 5800 12039 5808
rect 11494 5789 11527 5797
rect 11494 5772 11502 5789
rect 11519 5772 11527 5789
rect 11494 5764 11527 5772
rect 11861 5773 11894 5781
rect 11861 5756 11869 5773
rect 11886 5756 11894 5773
rect 11861 5748 11894 5756
rect 11911 5731 11938 5800
rect 12061 5731 12088 5854
rect 12522 6099 12580 6107
rect 12522 6082 12558 6099
rect 12575 6082 12580 6099
rect 12522 6065 12580 6082
rect 12522 6048 12558 6065
rect 12575 6048 12580 6065
rect 12522 6031 12580 6048
rect 12522 6014 12558 6031
rect 12575 6014 12580 6031
rect 12522 5997 12580 6014
rect 12522 5980 12558 5997
rect 12575 5980 12580 5997
rect 12522 5963 12580 5980
rect 12522 5946 12558 5963
rect 12575 5946 12580 5963
rect 12522 5929 12580 5946
rect 12522 5912 12558 5929
rect 12575 5912 12580 5929
rect 12522 5904 12580 5912
rect 12597 6099 12624 6122
rect 12597 6082 12602 6099
rect 12619 6082 12624 6099
rect 12597 6065 12624 6082
rect 12597 6048 12602 6065
rect 12619 6048 12624 6065
rect 12597 6031 12624 6048
rect 12597 6014 12602 6031
rect 12619 6014 12624 6031
rect 12597 5997 12624 6014
rect 12597 5980 12602 5997
rect 12619 5980 12624 5997
rect 12597 5963 12624 5980
rect 12597 5946 12602 5963
rect 12619 5946 12624 5963
rect 12597 5929 12624 5946
rect 12597 5912 12602 5929
rect 12619 5912 12624 5929
rect 12597 5904 12624 5912
rect 12641 6099 12699 6107
rect 12641 6082 12646 6099
rect 12663 6082 12699 6099
rect 12641 6065 12699 6082
rect 12641 6048 12646 6065
rect 12663 6048 12699 6065
rect 12641 6031 12699 6048
rect 12641 6014 12646 6031
rect 12663 6014 12699 6031
rect 12641 5997 12699 6014
rect 12641 5980 12646 5997
rect 12663 5980 12699 5997
rect 12641 5963 12699 5980
rect 12641 5946 12646 5963
rect 12663 5946 12699 5963
rect 12641 5929 12699 5946
rect 12641 5912 12646 5929
rect 12663 5912 12699 5929
rect 12641 5904 12699 5912
rect 12472 5827 12505 5835
rect 12472 5810 12480 5827
rect 12497 5810 12505 5827
rect 12472 5802 12505 5810
rect 12522 5817 12549 5904
rect 12571 5879 12604 5887
rect 12571 5862 12579 5879
rect 12596 5871 12604 5879
rect 12672 5871 12699 5904
rect 12596 5862 12699 5871
rect 12571 5854 12699 5862
rect 12617 5825 12650 5833
rect 12617 5817 12625 5825
rect 12522 5808 12625 5817
rect 12642 5808 12650 5825
rect 12522 5800 12650 5808
rect 12105 5789 12138 5797
rect 12105 5772 12113 5789
rect 12130 5772 12138 5789
rect 12105 5764 12138 5772
rect 12472 5773 12505 5781
rect 12472 5756 12480 5773
rect 12497 5756 12505 5773
rect 12472 5748 12505 5756
rect 12522 5731 12549 5800
rect 12672 5731 12699 5854
rect 12716 5789 12749 5797
rect 12716 5772 12724 5789
rect 12741 5772 12749 5789
rect 12716 5764 12749 5772
rect 9451 5723 9478 5731
rect 9451 5706 9456 5723
rect 9473 5706 9478 5723
rect 9451 5689 9478 5706
rect 9451 5672 9456 5689
rect 9473 5672 9478 5689
rect 9451 5655 9478 5672
rect 9451 5638 9456 5655
rect 9473 5638 9478 5655
rect 9451 5630 9478 5638
rect 9500 5723 9558 5731
rect 9500 5706 9536 5723
rect 9553 5706 9558 5723
rect 9500 5689 9558 5706
rect 9500 5672 9536 5689
rect 9553 5672 9558 5689
rect 9500 5655 9558 5672
rect 9500 5638 9536 5655
rect 9553 5638 9558 5655
rect 9500 5630 9558 5638
rect 9575 5723 9602 5731
rect 9575 5706 9580 5723
rect 9597 5706 9602 5723
rect 9575 5689 9602 5706
rect 9575 5672 9580 5689
rect 9597 5672 9602 5689
rect 9575 5655 9602 5672
rect 9575 5638 9580 5655
rect 9597 5638 9602 5655
rect 9575 5615 9602 5638
rect 9619 5723 9677 5731
rect 9619 5706 9624 5723
rect 9641 5706 9677 5723
rect 9619 5689 9677 5706
rect 9619 5672 9624 5689
rect 9641 5672 9677 5689
rect 9619 5655 9677 5672
rect 9619 5638 9624 5655
rect 9641 5638 9677 5655
rect 9619 5630 9677 5638
rect 9699 5723 9726 5731
rect 9699 5706 9704 5723
rect 9721 5706 9726 5723
rect 9699 5689 9726 5706
rect 9699 5672 9704 5689
rect 9721 5672 9726 5689
rect 9699 5655 9726 5672
rect 9699 5638 9704 5655
rect 9721 5638 9726 5655
rect 9699 5630 9726 5638
rect 10062 5723 10089 5731
rect 10062 5706 10067 5723
rect 10084 5706 10089 5723
rect 10062 5689 10089 5706
rect 10062 5672 10067 5689
rect 10084 5672 10089 5689
rect 10062 5655 10089 5672
rect 10062 5638 10067 5655
rect 10084 5638 10089 5655
rect 10062 5630 10089 5638
rect 10111 5723 10169 5731
rect 10111 5706 10147 5723
rect 10164 5706 10169 5723
rect 10111 5689 10169 5706
rect 10111 5672 10147 5689
rect 10164 5672 10169 5689
rect 10111 5655 10169 5672
rect 10111 5638 10147 5655
rect 10164 5638 10169 5655
rect 10111 5630 10169 5638
rect 10186 5723 10213 5731
rect 10186 5706 10191 5723
rect 10208 5706 10213 5723
rect 10186 5689 10213 5706
rect 10186 5672 10191 5689
rect 10208 5672 10213 5689
rect 10186 5655 10213 5672
rect 10186 5638 10191 5655
rect 10208 5638 10213 5655
rect 9575 5596 9579 5615
rect 9598 5596 9602 5615
rect 10186 5615 10213 5638
rect 10230 5723 10288 5731
rect 10230 5706 10235 5723
rect 10252 5706 10288 5723
rect 10230 5689 10288 5706
rect 10230 5672 10235 5689
rect 10252 5672 10288 5689
rect 10230 5655 10288 5672
rect 10230 5638 10235 5655
rect 10252 5638 10288 5655
rect 10230 5630 10288 5638
rect 10310 5723 10337 5731
rect 10310 5706 10315 5723
rect 10332 5706 10337 5723
rect 10310 5689 10337 5706
rect 10310 5672 10315 5689
rect 10332 5672 10337 5689
rect 10310 5655 10337 5672
rect 10310 5638 10315 5655
rect 10332 5638 10337 5655
rect 10310 5630 10337 5638
rect 10673 5723 10700 5731
rect 10673 5706 10678 5723
rect 10695 5706 10700 5723
rect 10673 5689 10700 5706
rect 10673 5672 10678 5689
rect 10695 5672 10700 5689
rect 10673 5655 10700 5672
rect 10673 5638 10678 5655
rect 10695 5638 10700 5655
rect 10673 5630 10700 5638
rect 10722 5723 10780 5731
rect 10722 5706 10758 5723
rect 10775 5706 10780 5723
rect 10722 5689 10780 5706
rect 10722 5672 10758 5689
rect 10775 5672 10780 5689
rect 10722 5655 10780 5672
rect 10722 5638 10758 5655
rect 10775 5638 10780 5655
rect 10722 5630 10780 5638
rect 10797 5723 10824 5731
rect 10797 5706 10802 5723
rect 10819 5706 10824 5723
rect 10797 5689 10824 5706
rect 10797 5672 10802 5689
rect 10819 5672 10824 5689
rect 10797 5655 10824 5672
rect 10797 5638 10802 5655
rect 10819 5638 10824 5655
rect 10186 5596 10190 5615
rect 10209 5596 10213 5615
rect 10797 5615 10824 5638
rect 10841 5723 10899 5731
rect 10841 5706 10846 5723
rect 10863 5706 10899 5723
rect 10841 5689 10899 5706
rect 10841 5672 10846 5689
rect 10863 5672 10899 5689
rect 10841 5655 10899 5672
rect 10841 5638 10846 5655
rect 10863 5638 10899 5655
rect 10841 5630 10899 5638
rect 10921 5723 10948 5731
rect 10921 5706 10926 5723
rect 10943 5706 10948 5723
rect 10921 5689 10948 5706
rect 10921 5672 10926 5689
rect 10943 5672 10948 5689
rect 10921 5655 10948 5672
rect 10921 5638 10926 5655
rect 10943 5638 10948 5655
rect 10921 5630 10948 5638
rect 11251 5723 11278 5731
rect 11251 5706 11256 5723
rect 11273 5706 11278 5723
rect 11251 5689 11278 5706
rect 11251 5672 11256 5689
rect 11273 5672 11278 5689
rect 11251 5655 11278 5672
rect 11251 5638 11256 5655
rect 11273 5638 11278 5655
rect 11251 5630 11278 5638
rect 11300 5723 11358 5731
rect 11300 5706 11336 5723
rect 11353 5706 11358 5723
rect 11300 5689 11358 5706
rect 11300 5672 11336 5689
rect 11353 5672 11358 5689
rect 11300 5655 11358 5672
rect 11300 5638 11336 5655
rect 11353 5638 11358 5655
rect 11300 5630 11358 5638
rect 11375 5723 11402 5731
rect 11375 5706 11380 5723
rect 11397 5706 11402 5723
rect 11375 5689 11402 5706
rect 11375 5672 11380 5689
rect 11397 5672 11402 5689
rect 11375 5655 11402 5672
rect 11375 5638 11380 5655
rect 11397 5638 11402 5655
rect 10797 5596 10801 5615
rect 10820 5596 10824 5615
rect 11375 5615 11402 5638
rect 11419 5723 11477 5731
rect 11419 5706 11424 5723
rect 11441 5706 11477 5723
rect 11419 5689 11477 5706
rect 11419 5672 11424 5689
rect 11441 5672 11477 5689
rect 11419 5655 11477 5672
rect 11419 5638 11424 5655
rect 11441 5638 11477 5655
rect 11419 5630 11477 5638
rect 11499 5723 11526 5731
rect 11499 5706 11504 5723
rect 11521 5706 11526 5723
rect 11499 5689 11526 5706
rect 11499 5672 11504 5689
rect 11521 5672 11526 5689
rect 11499 5655 11526 5672
rect 11499 5638 11504 5655
rect 11521 5638 11526 5655
rect 11499 5630 11526 5638
rect 11862 5723 11889 5731
rect 11862 5706 11867 5723
rect 11884 5706 11889 5723
rect 11862 5689 11889 5706
rect 11862 5672 11867 5689
rect 11884 5672 11889 5689
rect 11862 5655 11889 5672
rect 11862 5638 11867 5655
rect 11884 5638 11889 5655
rect 11862 5630 11889 5638
rect 11911 5723 11969 5731
rect 11911 5706 11947 5723
rect 11964 5706 11969 5723
rect 11911 5689 11969 5706
rect 11911 5672 11947 5689
rect 11964 5672 11969 5689
rect 11911 5655 11969 5672
rect 11911 5638 11947 5655
rect 11964 5638 11969 5655
rect 11911 5630 11969 5638
rect 11986 5723 12013 5731
rect 11986 5706 11991 5723
rect 12008 5706 12013 5723
rect 11986 5689 12013 5706
rect 11986 5672 11991 5689
rect 12008 5672 12013 5689
rect 11986 5655 12013 5672
rect 11986 5638 11991 5655
rect 12008 5638 12013 5655
rect 11375 5596 11379 5615
rect 11398 5596 11402 5615
rect 11986 5615 12013 5638
rect 12030 5723 12088 5731
rect 12030 5706 12035 5723
rect 12052 5706 12088 5723
rect 12030 5689 12088 5706
rect 12030 5672 12035 5689
rect 12052 5672 12088 5689
rect 12030 5655 12088 5672
rect 12030 5638 12035 5655
rect 12052 5638 12088 5655
rect 12030 5630 12088 5638
rect 12110 5723 12137 5731
rect 12110 5706 12115 5723
rect 12132 5706 12137 5723
rect 12110 5689 12137 5706
rect 12110 5672 12115 5689
rect 12132 5672 12137 5689
rect 12110 5655 12137 5672
rect 12110 5638 12115 5655
rect 12132 5638 12137 5655
rect 12110 5630 12137 5638
rect 12473 5723 12500 5731
rect 12473 5706 12478 5723
rect 12495 5706 12500 5723
rect 12473 5689 12500 5706
rect 12473 5672 12478 5689
rect 12495 5672 12500 5689
rect 12473 5655 12500 5672
rect 12473 5638 12478 5655
rect 12495 5638 12500 5655
rect 12473 5630 12500 5638
rect 12522 5723 12580 5731
rect 12522 5706 12558 5723
rect 12575 5706 12580 5723
rect 12522 5689 12580 5706
rect 12522 5672 12558 5689
rect 12575 5672 12580 5689
rect 12522 5655 12580 5672
rect 12522 5638 12558 5655
rect 12575 5638 12580 5655
rect 12522 5630 12580 5638
rect 12597 5723 12624 5731
rect 12597 5706 12602 5723
rect 12619 5706 12624 5723
rect 12597 5689 12624 5706
rect 12597 5672 12602 5689
rect 12619 5672 12624 5689
rect 12597 5655 12624 5672
rect 12597 5638 12602 5655
rect 12619 5638 12624 5655
rect 11986 5596 11990 5615
rect 12009 5596 12013 5615
rect 12597 5615 12624 5638
rect 12641 5723 12699 5731
rect 12641 5706 12646 5723
rect 12663 5706 12699 5723
rect 12641 5689 12699 5706
rect 12641 5672 12646 5689
rect 12663 5672 12699 5689
rect 12641 5655 12699 5672
rect 12641 5638 12646 5655
rect 12663 5638 12699 5655
rect 12641 5630 12699 5638
rect 12721 5723 12748 5731
rect 12721 5706 12726 5723
rect 12743 5706 12748 5723
rect 12721 5689 12748 5706
rect 12721 5672 12726 5689
rect 12743 5672 12748 5689
rect 12721 5655 12748 5672
rect 12721 5638 12726 5655
rect 12743 5638 12748 5655
rect 12721 5630 12748 5638
rect 12597 5596 12601 5615
rect 12620 5596 12624 5615
rect 9575 5472 9579 5491
rect 9598 5472 9602 5491
rect 9500 5449 9558 5457
rect 9500 5432 9536 5449
rect 9553 5432 9558 5449
rect 9500 5415 9558 5432
rect 9500 5398 9536 5415
rect 9553 5398 9558 5415
rect 9500 5381 9558 5398
rect 9500 5364 9536 5381
rect 9553 5364 9558 5381
rect 9500 5347 9558 5364
rect 9500 5330 9536 5347
rect 9553 5330 9558 5347
rect 9500 5313 9558 5330
rect 9500 5296 9536 5313
rect 9553 5296 9558 5313
rect 9500 5279 9558 5296
rect 9500 5262 9536 5279
rect 9553 5262 9558 5279
rect 9500 5254 9558 5262
rect 9575 5449 9602 5472
rect 10186 5472 10190 5491
rect 10209 5472 10213 5491
rect 9575 5432 9580 5449
rect 9597 5432 9602 5449
rect 9575 5415 9602 5432
rect 9575 5398 9580 5415
rect 9597 5398 9602 5415
rect 9575 5381 9602 5398
rect 9575 5364 9580 5381
rect 9597 5364 9602 5381
rect 9575 5347 9602 5364
rect 9575 5330 9580 5347
rect 9597 5330 9602 5347
rect 9575 5313 9602 5330
rect 9575 5296 9580 5313
rect 9597 5296 9602 5313
rect 9575 5279 9602 5296
rect 9575 5262 9580 5279
rect 9597 5262 9602 5279
rect 9575 5254 9602 5262
rect 9619 5449 9677 5457
rect 9619 5432 9624 5449
rect 9641 5432 9677 5449
rect 9619 5415 9677 5432
rect 9619 5398 9624 5415
rect 9641 5398 9677 5415
rect 9619 5381 9677 5398
rect 9619 5364 9624 5381
rect 9641 5364 9677 5381
rect 9619 5347 9677 5364
rect 9619 5330 9624 5347
rect 9641 5330 9677 5347
rect 9619 5313 9677 5330
rect 9619 5296 9624 5313
rect 9641 5296 9677 5313
rect 9619 5279 9677 5296
rect 9619 5262 9624 5279
rect 9641 5262 9677 5279
rect 9619 5254 9677 5262
rect 9450 5177 9483 5185
rect 9450 5160 9458 5177
rect 9475 5160 9483 5177
rect 9450 5152 9483 5160
rect 9500 5167 9527 5254
rect 9549 5229 9582 5237
rect 9549 5212 9557 5229
rect 9574 5221 9582 5229
rect 9650 5221 9677 5254
rect 9574 5212 9677 5221
rect 9549 5204 9677 5212
rect 9595 5175 9628 5183
rect 9595 5167 9603 5175
rect 9500 5158 9603 5167
rect 9620 5158 9628 5175
rect 9500 5150 9628 5158
rect 9450 5123 9483 5131
rect 9450 5106 9458 5123
rect 9475 5106 9483 5123
rect 9450 5098 9483 5106
rect 9500 5081 9527 5150
rect 9650 5081 9677 5204
rect 10111 5449 10169 5457
rect 10111 5432 10147 5449
rect 10164 5432 10169 5449
rect 10111 5415 10169 5432
rect 10111 5398 10147 5415
rect 10164 5398 10169 5415
rect 10111 5381 10169 5398
rect 10111 5364 10147 5381
rect 10164 5364 10169 5381
rect 10111 5347 10169 5364
rect 10111 5330 10147 5347
rect 10164 5330 10169 5347
rect 10111 5313 10169 5330
rect 10111 5296 10147 5313
rect 10164 5296 10169 5313
rect 10111 5279 10169 5296
rect 10111 5262 10147 5279
rect 10164 5262 10169 5279
rect 10111 5254 10169 5262
rect 10186 5449 10213 5472
rect 10797 5472 10801 5491
rect 10820 5472 10824 5491
rect 10186 5432 10191 5449
rect 10208 5432 10213 5449
rect 10186 5415 10213 5432
rect 10186 5398 10191 5415
rect 10208 5398 10213 5415
rect 10186 5381 10213 5398
rect 10186 5364 10191 5381
rect 10208 5364 10213 5381
rect 10186 5347 10213 5364
rect 10186 5330 10191 5347
rect 10208 5330 10213 5347
rect 10186 5313 10213 5330
rect 10186 5296 10191 5313
rect 10208 5296 10213 5313
rect 10186 5279 10213 5296
rect 10186 5262 10191 5279
rect 10208 5262 10213 5279
rect 10186 5254 10213 5262
rect 10230 5449 10288 5457
rect 10230 5432 10235 5449
rect 10252 5432 10288 5449
rect 10230 5415 10288 5432
rect 10230 5398 10235 5415
rect 10252 5398 10288 5415
rect 10230 5381 10288 5398
rect 10230 5364 10235 5381
rect 10252 5364 10288 5381
rect 10230 5347 10288 5364
rect 10230 5330 10235 5347
rect 10252 5330 10288 5347
rect 10230 5313 10288 5330
rect 10230 5296 10235 5313
rect 10252 5296 10288 5313
rect 10230 5279 10288 5296
rect 10230 5262 10235 5279
rect 10252 5262 10288 5279
rect 10230 5254 10288 5262
rect 10061 5177 10094 5185
rect 10061 5160 10069 5177
rect 10086 5160 10094 5177
rect 10061 5152 10094 5160
rect 10111 5167 10138 5254
rect 10160 5229 10193 5237
rect 10160 5212 10168 5229
rect 10185 5221 10193 5229
rect 10261 5221 10288 5254
rect 10185 5212 10288 5221
rect 10160 5204 10288 5212
rect 10206 5175 10239 5183
rect 10206 5167 10214 5175
rect 10111 5158 10214 5167
rect 10231 5158 10239 5175
rect 10111 5150 10239 5158
rect 9694 5139 9727 5147
rect 9694 5122 9702 5139
rect 9719 5122 9727 5139
rect 9694 5114 9727 5122
rect 10061 5123 10094 5131
rect 10061 5106 10069 5123
rect 10086 5106 10094 5123
rect 10061 5098 10094 5106
rect 10111 5081 10138 5150
rect 10261 5081 10288 5204
rect 10722 5449 10780 5457
rect 10722 5432 10758 5449
rect 10775 5432 10780 5449
rect 10722 5415 10780 5432
rect 10722 5398 10758 5415
rect 10775 5398 10780 5415
rect 10722 5381 10780 5398
rect 10722 5364 10758 5381
rect 10775 5364 10780 5381
rect 10722 5347 10780 5364
rect 10722 5330 10758 5347
rect 10775 5330 10780 5347
rect 10722 5313 10780 5330
rect 10722 5296 10758 5313
rect 10775 5296 10780 5313
rect 10722 5279 10780 5296
rect 10722 5262 10758 5279
rect 10775 5262 10780 5279
rect 10722 5254 10780 5262
rect 10797 5449 10824 5472
rect 11375 5472 11379 5491
rect 11398 5472 11402 5491
rect 10797 5432 10802 5449
rect 10819 5432 10824 5449
rect 10797 5415 10824 5432
rect 10797 5398 10802 5415
rect 10819 5398 10824 5415
rect 10797 5381 10824 5398
rect 10797 5364 10802 5381
rect 10819 5364 10824 5381
rect 10797 5347 10824 5364
rect 10797 5330 10802 5347
rect 10819 5330 10824 5347
rect 10797 5313 10824 5330
rect 10797 5296 10802 5313
rect 10819 5296 10824 5313
rect 10797 5279 10824 5296
rect 10797 5262 10802 5279
rect 10819 5262 10824 5279
rect 10797 5254 10824 5262
rect 10841 5449 10899 5457
rect 10841 5432 10846 5449
rect 10863 5432 10899 5449
rect 10841 5415 10899 5432
rect 10841 5398 10846 5415
rect 10863 5398 10899 5415
rect 10841 5381 10899 5398
rect 10841 5364 10846 5381
rect 10863 5364 10899 5381
rect 10841 5347 10899 5364
rect 10841 5330 10846 5347
rect 10863 5330 10899 5347
rect 10841 5313 10899 5330
rect 10841 5296 10846 5313
rect 10863 5296 10899 5313
rect 10841 5279 10899 5296
rect 10841 5262 10846 5279
rect 10863 5262 10899 5279
rect 10841 5254 10899 5262
rect 10672 5177 10705 5185
rect 10672 5160 10680 5177
rect 10697 5160 10705 5177
rect 10672 5152 10705 5160
rect 10722 5167 10749 5254
rect 10771 5229 10804 5237
rect 10771 5212 10779 5229
rect 10796 5221 10804 5229
rect 10872 5221 10899 5254
rect 10796 5212 10899 5221
rect 10771 5204 10899 5212
rect 10817 5175 10850 5183
rect 10817 5167 10825 5175
rect 10722 5158 10825 5167
rect 10842 5158 10850 5175
rect 10722 5150 10850 5158
rect 10305 5139 10338 5147
rect 10305 5122 10313 5139
rect 10330 5122 10338 5139
rect 10305 5114 10338 5122
rect 10672 5123 10705 5131
rect 10672 5106 10680 5123
rect 10697 5106 10705 5123
rect 10672 5098 10705 5106
rect 10722 5081 10749 5150
rect 10872 5081 10899 5204
rect 11300 5449 11358 5457
rect 11300 5432 11336 5449
rect 11353 5432 11358 5449
rect 11300 5415 11358 5432
rect 11300 5398 11336 5415
rect 11353 5398 11358 5415
rect 11300 5381 11358 5398
rect 11300 5364 11336 5381
rect 11353 5364 11358 5381
rect 11300 5347 11358 5364
rect 11300 5330 11336 5347
rect 11353 5330 11358 5347
rect 11300 5313 11358 5330
rect 11300 5296 11336 5313
rect 11353 5296 11358 5313
rect 11300 5279 11358 5296
rect 11300 5262 11336 5279
rect 11353 5262 11358 5279
rect 11300 5254 11358 5262
rect 11375 5449 11402 5472
rect 11986 5472 11990 5491
rect 12009 5472 12013 5491
rect 11375 5432 11380 5449
rect 11397 5432 11402 5449
rect 11375 5415 11402 5432
rect 11375 5398 11380 5415
rect 11397 5398 11402 5415
rect 11375 5381 11402 5398
rect 11375 5364 11380 5381
rect 11397 5364 11402 5381
rect 11375 5347 11402 5364
rect 11375 5330 11380 5347
rect 11397 5330 11402 5347
rect 11375 5313 11402 5330
rect 11375 5296 11380 5313
rect 11397 5296 11402 5313
rect 11375 5279 11402 5296
rect 11375 5262 11380 5279
rect 11397 5262 11402 5279
rect 11375 5254 11402 5262
rect 11419 5449 11477 5457
rect 11419 5432 11424 5449
rect 11441 5432 11477 5449
rect 11419 5415 11477 5432
rect 11419 5398 11424 5415
rect 11441 5398 11477 5415
rect 11419 5381 11477 5398
rect 11419 5364 11424 5381
rect 11441 5364 11477 5381
rect 11419 5347 11477 5364
rect 11419 5330 11424 5347
rect 11441 5330 11477 5347
rect 11419 5313 11477 5330
rect 11419 5296 11424 5313
rect 11441 5296 11477 5313
rect 11419 5279 11477 5296
rect 11419 5262 11424 5279
rect 11441 5262 11477 5279
rect 11419 5254 11477 5262
rect 11250 5177 11283 5185
rect 11250 5160 11258 5177
rect 11275 5160 11283 5177
rect 11250 5152 11283 5160
rect 11300 5167 11327 5254
rect 11349 5229 11382 5237
rect 11349 5212 11357 5229
rect 11374 5221 11382 5229
rect 11450 5221 11477 5254
rect 11374 5212 11477 5221
rect 11349 5204 11477 5212
rect 11395 5175 11428 5183
rect 11395 5167 11403 5175
rect 11300 5158 11403 5167
rect 11420 5158 11428 5175
rect 11300 5150 11428 5158
rect 10916 5139 10949 5147
rect 10916 5122 10924 5139
rect 10941 5122 10949 5139
rect 10916 5114 10949 5122
rect 11250 5123 11283 5131
rect 11250 5106 11258 5123
rect 11275 5106 11283 5123
rect 11250 5098 11283 5106
rect 11300 5081 11327 5150
rect 11450 5081 11477 5204
rect 11911 5449 11969 5457
rect 11911 5432 11947 5449
rect 11964 5432 11969 5449
rect 11911 5415 11969 5432
rect 11911 5398 11947 5415
rect 11964 5398 11969 5415
rect 11911 5381 11969 5398
rect 11911 5364 11947 5381
rect 11964 5364 11969 5381
rect 11911 5347 11969 5364
rect 11911 5330 11947 5347
rect 11964 5330 11969 5347
rect 11911 5313 11969 5330
rect 11911 5296 11947 5313
rect 11964 5296 11969 5313
rect 11911 5279 11969 5296
rect 11911 5262 11947 5279
rect 11964 5262 11969 5279
rect 11911 5254 11969 5262
rect 11986 5449 12013 5472
rect 12597 5472 12601 5491
rect 12620 5472 12624 5491
rect 11986 5432 11991 5449
rect 12008 5432 12013 5449
rect 11986 5415 12013 5432
rect 11986 5398 11991 5415
rect 12008 5398 12013 5415
rect 11986 5381 12013 5398
rect 11986 5364 11991 5381
rect 12008 5364 12013 5381
rect 11986 5347 12013 5364
rect 11986 5330 11991 5347
rect 12008 5330 12013 5347
rect 11986 5313 12013 5330
rect 11986 5296 11991 5313
rect 12008 5296 12013 5313
rect 11986 5279 12013 5296
rect 11986 5262 11991 5279
rect 12008 5262 12013 5279
rect 11986 5254 12013 5262
rect 12030 5449 12088 5457
rect 12030 5432 12035 5449
rect 12052 5432 12088 5449
rect 12030 5415 12088 5432
rect 12030 5398 12035 5415
rect 12052 5398 12088 5415
rect 12030 5381 12088 5398
rect 12030 5364 12035 5381
rect 12052 5364 12088 5381
rect 12030 5347 12088 5364
rect 12030 5330 12035 5347
rect 12052 5330 12088 5347
rect 12030 5313 12088 5330
rect 12030 5296 12035 5313
rect 12052 5296 12088 5313
rect 12030 5279 12088 5296
rect 12030 5262 12035 5279
rect 12052 5262 12088 5279
rect 12030 5254 12088 5262
rect 11861 5177 11894 5185
rect 11861 5160 11869 5177
rect 11886 5160 11894 5177
rect 11861 5152 11894 5160
rect 11911 5167 11938 5254
rect 11960 5229 11993 5237
rect 11960 5212 11968 5229
rect 11985 5221 11993 5229
rect 12061 5221 12088 5254
rect 11985 5212 12088 5221
rect 11960 5204 12088 5212
rect 12006 5175 12039 5183
rect 12006 5167 12014 5175
rect 11911 5158 12014 5167
rect 12031 5158 12039 5175
rect 11911 5150 12039 5158
rect 11494 5139 11527 5147
rect 11494 5122 11502 5139
rect 11519 5122 11527 5139
rect 11494 5114 11527 5122
rect 11861 5123 11894 5131
rect 11861 5106 11869 5123
rect 11886 5106 11894 5123
rect 11861 5098 11894 5106
rect 11911 5081 11938 5150
rect 12061 5081 12088 5204
rect 12522 5449 12580 5457
rect 12522 5432 12558 5449
rect 12575 5432 12580 5449
rect 12522 5415 12580 5432
rect 12522 5398 12558 5415
rect 12575 5398 12580 5415
rect 12522 5381 12580 5398
rect 12522 5364 12558 5381
rect 12575 5364 12580 5381
rect 12522 5347 12580 5364
rect 12522 5330 12558 5347
rect 12575 5330 12580 5347
rect 12522 5313 12580 5330
rect 12522 5296 12558 5313
rect 12575 5296 12580 5313
rect 12522 5279 12580 5296
rect 12522 5262 12558 5279
rect 12575 5262 12580 5279
rect 12522 5254 12580 5262
rect 12597 5449 12624 5472
rect 12597 5432 12602 5449
rect 12619 5432 12624 5449
rect 12597 5415 12624 5432
rect 12597 5398 12602 5415
rect 12619 5398 12624 5415
rect 12597 5381 12624 5398
rect 12597 5364 12602 5381
rect 12619 5364 12624 5381
rect 12597 5347 12624 5364
rect 12597 5330 12602 5347
rect 12619 5330 12624 5347
rect 12597 5313 12624 5330
rect 12597 5296 12602 5313
rect 12619 5296 12624 5313
rect 12597 5279 12624 5296
rect 12597 5262 12602 5279
rect 12619 5262 12624 5279
rect 12597 5254 12624 5262
rect 12641 5449 12699 5457
rect 12641 5432 12646 5449
rect 12663 5432 12699 5449
rect 12641 5415 12699 5432
rect 12641 5398 12646 5415
rect 12663 5398 12699 5415
rect 12641 5381 12699 5398
rect 12641 5364 12646 5381
rect 12663 5364 12699 5381
rect 12641 5347 12699 5364
rect 12641 5330 12646 5347
rect 12663 5330 12699 5347
rect 12641 5313 12699 5330
rect 12641 5296 12646 5313
rect 12663 5296 12699 5313
rect 12641 5279 12699 5296
rect 12641 5262 12646 5279
rect 12663 5262 12699 5279
rect 12641 5254 12699 5262
rect 12472 5177 12505 5185
rect 12472 5160 12480 5177
rect 12497 5160 12505 5177
rect 12472 5152 12505 5160
rect 12522 5167 12549 5254
rect 12571 5229 12604 5237
rect 12571 5212 12579 5229
rect 12596 5221 12604 5229
rect 12672 5221 12699 5254
rect 12596 5212 12699 5221
rect 12571 5204 12699 5212
rect 12617 5175 12650 5183
rect 12617 5167 12625 5175
rect 12522 5158 12625 5167
rect 12642 5158 12650 5175
rect 12522 5150 12650 5158
rect 12105 5139 12138 5147
rect 12105 5122 12113 5139
rect 12130 5122 12138 5139
rect 12105 5114 12138 5122
rect 12472 5123 12505 5131
rect 12472 5106 12480 5123
rect 12497 5106 12505 5123
rect 12472 5098 12505 5106
rect 12522 5081 12549 5150
rect 12672 5081 12699 5204
rect 12716 5139 12749 5147
rect 12716 5122 12724 5139
rect 12741 5122 12749 5139
rect 12716 5114 12749 5122
rect 9451 5073 9478 5081
rect 9451 5056 9456 5073
rect 9473 5056 9478 5073
rect 9451 5039 9478 5056
rect 9451 5022 9456 5039
rect 9473 5022 9478 5039
rect 9451 5005 9478 5022
rect 9451 4988 9456 5005
rect 9473 4988 9478 5005
rect 9451 4980 9478 4988
rect 9500 5073 9558 5081
rect 9500 5056 9536 5073
rect 9553 5056 9558 5073
rect 9500 5039 9558 5056
rect 9500 5022 9536 5039
rect 9553 5022 9558 5039
rect 9500 5005 9558 5022
rect 9500 4988 9536 5005
rect 9553 4988 9558 5005
rect 9500 4980 9558 4988
rect 9575 5073 9602 5081
rect 9575 5056 9580 5073
rect 9597 5056 9602 5073
rect 9575 5039 9602 5056
rect 9575 5022 9580 5039
rect 9597 5022 9602 5039
rect 9575 5005 9602 5022
rect 9575 4988 9580 5005
rect 9597 4988 9602 5005
rect 9575 4965 9602 4988
rect 9619 5073 9677 5081
rect 9619 5056 9624 5073
rect 9641 5056 9677 5073
rect 9619 5039 9677 5056
rect 9619 5022 9624 5039
rect 9641 5022 9677 5039
rect 9619 5005 9677 5022
rect 9619 4988 9624 5005
rect 9641 4988 9677 5005
rect 9619 4980 9677 4988
rect 9699 5073 9726 5081
rect 9699 5056 9704 5073
rect 9721 5056 9726 5073
rect 9699 5039 9726 5056
rect 9699 5022 9704 5039
rect 9721 5022 9726 5039
rect 9699 5005 9726 5022
rect 9699 4988 9704 5005
rect 9721 4988 9726 5005
rect 9699 4980 9726 4988
rect 10062 5073 10089 5081
rect 10062 5056 10067 5073
rect 10084 5056 10089 5073
rect 10062 5039 10089 5056
rect 10062 5022 10067 5039
rect 10084 5022 10089 5039
rect 10062 5005 10089 5022
rect 10062 4988 10067 5005
rect 10084 4988 10089 5005
rect 10062 4980 10089 4988
rect 10111 5073 10169 5081
rect 10111 5056 10147 5073
rect 10164 5056 10169 5073
rect 10111 5039 10169 5056
rect 10111 5022 10147 5039
rect 10164 5022 10169 5039
rect 10111 5005 10169 5022
rect 10111 4988 10147 5005
rect 10164 4988 10169 5005
rect 10111 4980 10169 4988
rect 10186 5073 10213 5081
rect 10186 5056 10191 5073
rect 10208 5056 10213 5073
rect 10186 5039 10213 5056
rect 10186 5022 10191 5039
rect 10208 5022 10213 5039
rect 10186 5005 10213 5022
rect 10186 4988 10191 5005
rect 10208 4988 10213 5005
rect 9575 4946 9579 4965
rect 9598 4946 9602 4965
rect 10186 4965 10213 4988
rect 10230 5073 10288 5081
rect 10230 5056 10235 5073
rect 10252 5056 10288 5073
rect 10230 5039 10288 5056
rect 10230 5022 10235 5039
rect 10252 5022 10288 5039
rect 10230 5005 10288 5022
rect 10230 4988 10235 5005
rect 10252 4988 10288 5005
rect 10230 4980 10288 4988
rect 10310 5073 10337 5081
rect 10310 5056 10315 5073
rect 10332 5056 10337 5073
rect 10310 5039 10337 5056
rect 10310 5022 10315 5039
rect 10332 5022 10337 5039
rect 10310 5005 10337 5022
rect 10310 4988 10315 5005
rect 10332 4988 10337 5005
rect 10310 4980 10337 4988
rect 10673 5073 10700 5081
rect 10673 5056 10678 5073
rect 10695 5056 10700 5073
rect 10673 5039 10700 5056
rect 10673 5022 10678 5039
rect 10695 5022 10700 5039
rect 10673 5005 10700 5022
rect 10673 4988 10678 5005
rect 10695 4988 10700 5005
rect 10673 4980 10700 4988
rect 10722 5073 10780 5081
rect 10722 5056 10758 5073
rect 10775 5056 10780 5073
rect 10722 5039 10780 5056
rect 10722 5022 10758 5039
rect 10775 5022 10780 5039
rect 10722 5005 10780 5022
rect 10722 4988 10758 5005
rect 10775 4988 10780 5005
rect 10722 4980 10780 4988
rect 10797 5073 10824 5081
rect 10797 5056 10802 5073
rect 10819 5056 10824 5073
rect 10797 5039 10824 5056
rect 10797 5022 10802 5039
rect 10819 5022 10824 5039
rect 10797 5005 10824 5022
rect 10797 4988 10802 5005
rect 10819 4988 10824 5005
rect 10186 4946 10190 4965
rect 10209 4946 10213 4965
rect 10797 4965 10824 4988
rect 10841 5073 10899 5081
rect 10841 5056 10846 5073
rect 10863 5056 10899 5073
rect 10841 5039 10899 5056
rect 10841 5022 10846 5039
rect 10863 5022 10899 5039
rect 10841 5005 10899 5022
rect 10841 4988 10846 5005
rect 10863 4988 10899 5005
rect 10841 4980 10899 4988
rect 10921 5073 10948 5081
rect 10921 5056 10926 5073
rect 10943 5056 10948 5073
rect 10921 5039 10948 5056
rect 10921 5022 10926 5039
rect 10943 5022 10948 5039
rect 10921 5005 10948 5022
rect 10921 4988 10926 5005
rect 10943 4988 10948 5005
rect 10921 4980 10948 4988
rect 11251 5073 11278 5081
rect 11251 5056 11256 5073
rect 11273 5056 11278 5073
rect 11251 5039 11278 5056
rect 11251 5022 11256 5039
rect 11273 5022 11278 5039
rect 11251 5005 11278 5022
rect 11251 4988 11256 5005
rect 11273 4988 11278 5005
rect 11251 4980 11278 4988
rect 11300 5073 11358 5081
rect 11300 5056 11336 5073
rect 11353 5056 11358 5073
rect 11300 5039 11358 5056
rect 11300 5022 11336 5039
rect 11353 5022 11358 5039
rect 11300 5005 11358 5022
rect 11300 4988 11336 5005
rect 11353 4988 11358 5005
rect 11300 4980 11358 4988
rect 11375 5073 11402 5081
rect 11375 5056 11380 5073
rect 11397 5056 11402 5073
rect 11375 5039 11402 5056
rect 11375 5022 11380 5039
rect 11397 5022 11402 5039
rect 11375 5005 11402 5022
rect 11375 4988 11380 5005
rect 11397 4988 11402 5005
rect 10797 4946 10801 4965
rect 10820 4946 10824 4965
rect 11375 4965 11402 4988
rect 11419 5073 11477 5081
rect 11419 5056 11424 5073
rect 11441 5056 11477 5073
rect 11419 5039 11477 5056
rect 11419 5022 11424 5039
rect 11441 5022 11477 5039
rect 11419 5005 11477 5022
rect 11419 4988 11424 5005
rect 11441 4988 11477 5005
rect 11419 4980 11477 4988
rect 11499 5073 11526 5081
rect 11499 5056 11504 5073
rect 11521 5056 11526 5073
rect 11499 5039 11526 5056
rect 11499 5022 11504 5039
rect 11521 5022 11526 5039
rect 11499 5005 11526 5022
rect 11499 4988 11504 5005
rect 11521 4988 11526 5005
rect 11499 4980 11526 4988
rect 11862 5073 11889 5081
rect 11862 5056 11867 5073
rect 11884 5056 11889 5073
rect 11862 5039 11889 5056
rect 11862 5022 11867 5039
rect 11884 5022 11889 5039
rect 11862 5005 11889 5022
rect 11862 4988 11867 5005
rect 11884 4988 11889 5005
rect 11862 4980 11889 4988
rect 11911 5073 11969 5081
rect 11911 5056 11947 5073
rect 11964 5056 11969 5073
rect 11911 5039 11969 5056
rect 11911 5022 11947 5039
rect 11964 5022 11969 5039
rect 11911 5005 11969 5022
rect 11911 4988 11947 5005
rect 11964 4988 11969 5005
rect 11911 4980 11969 4988
rect 11986 5073 12013 5081
rect 11986 5056 11991 5073
rect 12008 5056 12013 5073
rect 11986 5039 12013 5056
rect 11986 5022 11991 5039
rect 12008 5022 12013 5039
rect 11986 5005 12013 5022
rect 11986 4988 11991 5005
rect 12008 4988 12013 5005
rect 11375 4946 11379 4965
rect 11398 4946 11402 4965
rect 11986 4965 12013 4988
rect 12030 5073 12088 5081
rect 12030 5056 12035 5073
rect 12052 5056 12088 5073
rect 12030 5039 12088 5056
rect 12030 5022 12035 5039
rect 12052 5022 12088 5039
rect 12030 5005 12088 5022
rect 12030 4988 12035 5005
rect 12052 4988 12088 5005
rect 12030 4980 12088 4988
rect 12110 5073 12137 5081
rect 12110 5056 12115 5073
rect 12132 5056 12137 5073
rect 12110 5039 12137 5056
rect 12110 5022 12115 5039
rect 12132 5022 12137 5039
rect 12110 5005 12137 5022
rect 12110 4988 12115 5005
rect 12132 4988 12137 5005
rect 12110 4980 12137 4988
rect 12473 5073 12500 5081
rect 12473 5056 12478 5073
rect 12495 5056 12500 5073
rect 12473 5039 12500 5056
rect 12473 5022 12478 5039
rect 12495 5022 12500 5039
rect 12473 5005 12500 5022
rect 12473 4988 12478 5005
rect 12495 4988 12500 5005
rect 12473 4980 12500 4988
rect 12522 5073 12580 5081
rect 12522 5056 12558 5073
rect 12575 5056 12580 5073
rect 12522 5039 12580 5056
rect 12522 5022 12558 5039
rect 12575 5022 12580 5039
rect 12522 5005 12580 5022
rect 12522 4988 12558 5005
rect 12575 4988 12580 5005
rect 12522 4980 12580 4988
rect 12597 5073 12624 5081
rect 12597 5056 12602 5073
rect 12619 5056 12624 5073
rect 12597 5039 12624 5056
rect 12597 5022 12602 5039
rect 12619 5022 12624 5039
rect 12597 5005 12624 5022
rect 12597 4988 12602 5005
rect 12619 4988 12624 5005
rect 11986 4946 11990 4965
rect 12009 4946 12013 4965
rect 12597 4965 12624 4988
rect 12641 5073 12699 5081
rect 12641 5056 12646 5073
rect 12663 5056 12699 5073
rect 12641 5039 12699 5056
rect 12641 5022 12646 5039
rect 12663 5022 12699 5039
rect 12641 5005 12699 5022
rect 12641 4988 12646 5005
rect 12663 4988 12699 5005
rect 12641 4980 12699 4988
rect 12721 5073 12748 5081
rect 12721 5056 12726 5073
rect 12743 5056 12748 5073
rect 12721 5039 12748 5056
rect 12721 5022 12726 5039
rect 12743 5022 12748 5039
rect 12721 5005 12748 5022
rect 12721 4988 12726 5005
rect 12743 4988 12748 5005
rect 12721 4980 12748 4988
rect 12597 4946 12601 4965
rect 12620 4946 12624 4965
rect 9575 4832 9579 4851
rect 9598 4832 9602 4851
rect 9500 4809 9558 4817
rect 9500 4792 9536 4809
rect 9553 4792 9558 4809
rect 9500 4775 9558 4792
rect 9500 4758 9536 4775
rect 9553 4758 9558 4775
rect 9500 4741 9558 4758
rect 9500 4724 9536 4741
rect 9553 4724 9558 4741
rect 9500 4707 9558 4724
rect 9500 4690 9536 4707
rect 9553 4690 9558 4707
rect 9500 4673 9558 4690
rect 9500 4656 9536 4673
rect 9553 4656 9558 4673
rect 9500 4639 9558 4656
rect 9500 4622 9536 4639
rect 9553 4622 9558 4639
rect 9500 4614 9558 4622
rect 9575 4809 9602 4832
rect 10186 4832 10190 4851
rect 10209 4832 10213 4851
rect 9575 4792 9580 4809
rect 9597 4792 9602 4809
rect 9575 4775 9602 4792
rect 9575 4758 9580 4775
rect 9597 4758 9602 4775
rect 9575 4741 9602 4758
rect 9575 4724 9580 4741
rect 9597 4724 9602 4741
rect 9575 4707 9602 4724
rect 9575 4690 9580 4707
rect 9597 4690 9602 4707
rect 9575 4673 9602 4690
rect 9575 4656 9580 4673
rect 9597 4656 9602 4673
rect 9575 4639 9602 4656
rect 9575 4622 9580 4639
rect 9597 4622 9602 4639
rect 9575 4614 9602 4622
rect 9619 4809 9677 4817
rect 9619 4792 9624 4809
rect 9641 4792 9677 4809
rect 9619 4775 9677 4792
rect 9619 4758 9624 4775
rect 9641 4758 9677 4775
rect 9619 4741 9677 4758
rect 9619 4724 9624 4741
rect 9641 4724 9677 4741
rect 9619 4707 9677 4724
rect 9619 4690 9624 4707
rect 9641 4690 9677 4707
rect 9619 4673 9677 4690
rect 9619 4656 9624 4673
rect 9641 4656 9677 4673
rect 9619 4639 9677 4656
rect 9619 4622 9624 4639
rect 9641 4622 9677 4639
rect 9619 4614 9677 4622
rect 9450 4537 9483 4545
rect 9450 4520 9458 4537
rect 9475 4520 9483 4537
rect 9450 4512 9483 4520
rect 9500 4527 9527 4614
rect 9549 4589 9582 4597
rect 9549 4572 9557 4589
rect 9574 4581 9582 4589
rect 9650 4581 9677 4614
rect 9574 4572 9677 4581
rect 9549 4564 9677 4572
rect 9595 4535 9628 4543
rect 9595 4527 9603 4535
rect 9500 4518 9603 4527
rect 9620 4518 9628 4535
rect 9500 4510 9628 4518
rect 9450 4483 9483 4491
rect 9450 4466 9458 4483
rect 9475 4466 9483 4483
rect 9450 4458 9483 4466
rect 9500 4441 9527 4510
rect 9650 4441 9677 4564
rect 10111 4809 10169 4817
rect 10111 4792 10147 4809
rect 10164 4792 10169 4809
rect 10111 4775 10169 4792
rect 10111 4758 10147 4775
rect 10164 4758 10169 4775
rect 10111 4741 10169 4758
rect 10111 4724 10147 4741
rect 10164 4724 10169 4741
rect 10111 4707 10169 4724
rect 10111 4690 10147 4707
rect 10164 4690 10169 4707
rect 10111 4673 10169 4690
rect 10111 4656 10147 4673
rect 10164 4656 10169 4673
rect 10111 4639 10169 4656
rect 10111 4622 10147 4639
rect 10164 4622 10169 4639
rect 10111 4614 10169 4622
rect 10186 4809 10213 4832
rect 10797 4832 10801 4851
rect 10820 4832 10824 4851
rect 10186 4792 10191 4809
rect 10208 4792 10213 4809
rect 10186 4775 10213 4792
rect 10186 4758 10191 4775
rect 10208 4758 10213 4775
rect 10186 4741 10213 4758
rect 10186 4724 10191 4741
rect 10208 4724 10213 4741
rect 10186 4707 10213 4724
rect 10186 4690 10191 4707
rect 10208 4690 10213 4707
rect 10186 4673 10213 4690
rect 10186 4656 10191 4673
rect 10208 4656 10213 4673
rect 10186 4639 10213 4656
rect 10186 4622 10191 4639
rect 10208 4622 10213 4639
rect 10186 4614 10213 4622
rect 10230 4809 10288 4817
rect 10230 4792 10235 4809
rect 10252 4792 10288 4809
rect 10230 4775 10288 4792
rect 10230 4758 10235 4775
rect 10252 4758 10288 4775
rect 10230 4741 10288 4758
rect 10230 4724 10235 4741
rect 10252 4724 10288 4741
rect 10230 4707 10288 4724
rect 10230 4690 10235 4707
rect 10252 4690 10288 4707
rect 10230 4673 10288 4690
rect 10230 4656 10235 4673
rect 10252 4656 10288 4673
rect 10230 4639 10288 4656
rect 10230 4622 10235 4639
rect 10252 4622 10288 4639
rect 10230 4614 10288 4622
rect 10061 4537 10094 4545
rect 10061 4520 10069 4537
rect 10086 4520 10094 4537
rect 10061 4512 10094 4520
rect 10111 4527 10138 4614
rect 10160 4589 10193 4597
rect 10160 4572 10168 4589
rect 10185 4581 10193 4589
rect 10261 4581 10288 4614
rect 10185 4572 10288 4581
rect 10160 4564 10288 4572
rect 10206 4535 10239 4543
rect 10206 4527 10214 4535
rect 10111 4518 10214 4527
rect 10231 4518 10239 4535
rect 10111 4510 10239 4518
rect 9694 4499 9727 4507
rect 9694 4482 9702 4499
rect 9719 4482 9727 4499
rect 9694 4474 9727 4482
rect 10061 4483 10094 4491
rect 10061 4466 10069 4483
rect 10086 4466 10094 4483
rect 10061 4458 10094 4466
rect 10111 4441 10138 4510
rect 10261 4441 10288 4564
rect 10722 4809 10780 4817
rect 10722 4792 10758 4809
rect 10775 4792 10780 4809
rect 10722 4775 10780 4792
rect 10722 4758 10758 4775
rect 10775 4758 10780 4775
rect 10722 4741 10780 4758
rect 10722 4724 10758 4741
rect 10775 4724 10780 4741
rect 10722 4707 10780 4724
rect 10722 4690 10758 4707
rect 10775 4690 10780 4707
rect 10722 4673 10780 4690
rect 10722 4656 10758 4673
rect 10775 4656 10780 4673
rect 10722 4639 10780 4656
rect 10722 4622 10758 4639
rect 10775 4622 10780 4639
rect 10722 4614 10780 4622
rect 10797 4809 10824 4832
rect 11375 4832 11379 4851
rect 11398 4832 11402 4851
rect 10797 4792 10802 4809
rect 10819 4792 10824 4809
rect 10797 4775 10824 4792
rect 10797 4758 10802 4775
rect 10819 4758 10824 4775
rect 10797 4741 10824 4758
rect 10797 4724 10802 4741
rect 10819 4724 10824 4741
rect 10797 4707 10824 4724
rect 10797 4690 10802 4707
rect 10819 4690 10824 4707
rect 10797 4673 10824 4690
rect 10797 4656 10802 4673
rect 10819 4656 10824 4673
rect 10797 4639 10824 4656
rect 10797 4622 10802 4639
rect 10819 4622 10824 4639
rect 10797 4614 10824 4622
rect 10841 4809 10899 4817
rect 10841 4792 10846 4809
rect 10863 4792 10899 4809
rect 10841 4775 10899 4792
rect 10841 4758 10846 4775
rect 10863 4758 10899 4775
rect 10841 4741 10899 4758
rect 10841 4724 10846 4741
rect 10863 4724 10899 4741
rect 10841 4707 10899 4724
rect 10841 4690 10846 4707
rect 10863 4690 10899 4707
rect 10841 4673 10899 4690
rect 10841 4656 10846 4673
rect 10863 4656 10899 4673
rect 10841 4639 10899 4656
rect 10841 4622 10846 4639
rect 10863 4622 10899 4639
rect 10841 4614 10899 4622
rect 10672 4537 10705 4545
rect 10672 4520 10680 4537
rect 10697 4520 10705 4537
rect 10672 4512 10705 4520
rect 10722 4527 10749 4614
rect 10771 4589 10804 4597
rect 10771 4572 10779 4589
rect 10796 4581 10804 4589
rect 10872 4581 10899 4614
rect 10796 4572 10899 4581
rect 10771 4564 10899 4572
rect 10817 4535 10850 4543
rect 10817 4527 10825 4535
rect 10722 4518 10825 4527
rect 10842 4518 10850 4535
rect 10722 4510 10850 4518
rect 10305 4499 10338 4507
rect 10305 4482 10313 4499
rect 10330 4482 10338 4499
rect 10305 4474 10338 4482
rect 10672 4483 10705 4491
rect 10672 4466 10680 4483
rect 10697 4466 10705 4483
rect 10672 4458 10705 4466
rect 10722 4441 10749 4510
rect 10872 4441 10899 4564
rect 11300 4809 11358 4817
rect 11300 4792 11336 4809
rect 11353 4792 11358 4809
rect 11300 4775 11358 4792
rect 11300 4758 11336 4775
rect 11353 4758 11358 4775
rect 11300 4741 11358 4758
rect 11300 4724 11336 4741
rect 11353 4724 11358 4741
rect 11300 4707 11358 4724
rect 11300 4690 11336 4707
rect 11353 4690 11358 4707
rect 11300 4673 11358 4690
rect 11300 4656 11336 4673
rect 11353 4656 11358 4673
rect 11300 4639 11358 4656
rect 11300 4622 11336 4639
rect 11353 4622 11358 4639
rect 11300 4614 11358 4622
rect 11375 4809 11402 4832
rect 11986 4832 11990 4851
rect 12009 4832 12013 4851
rect 11375 4792 11380 4809
rect 11397 4792 11402 4809
rect 11375 4775 11402 4792
rect 11375 4758 11380 4775
rect 11397 4758 11402 4775
rect 11375 4741 11402 4758
rect 11375 4724 11380 4741
rect 11397 4724 11402 4741
rect 11375 4707 11402 4724
rect 11375 4690 11380 4707
rect 11397 4690 11402 4707
rect 11375 4673 11402 4690
rect 11375 4656 11380 4673
rect 11397 4656 11402 4673
rect 11375 4639 11402 4656
rect 11375 4622 11380 4639
rect 11397 4622 11402 4639
rect 11375 4614 11402 4622
rect 11419 4809 11477 4817
rect 11419 4792 11424 4809
rect 11441 4792 11477 4809
rect 11419 4775 11477 4792
rect 11419 4758 11424 4775
rect 11441 4758 11477 4775
rect 11419 4741 11477 4758
rect 11419 4724 11424 4741
rect 11441 4724 11477 4741
rect 11419 4707 11477 4724
rect 11419 4690 11424 4707
rect 11441 4690 11477 4707
rect 11419 4673 11477 4690
rect 11419 4656 11424 4673
rect 11441 4656 11477 4673
rect 11419 4639 11477 4656
rect 11419 4622 11424 4639
rect 11441 4622 11477 4639
rect 11419 4614 11477 4622
rect 11250 4537 11283 4545
rect 11250 4520 11258 4537
rect 11275 4520 11283 4537
rect 11250 4512 11283 4520
rect 11300 4527 11327 4614
rect 11349 4589 11382 4597
rect 11349 4572 11357 4589
rect 11374 4581 11382 4589
rect 11450 4581 11477 4614
rect 11374 4572 11477 4581
rect 11349 4564 11477 4572
rect 11395 4535 11428 4543
rect 11395 4527 11403 4535
rect 11300 4518 11403 4527
rect 11420 4518 11428 4535
rect 11300 4510 11428 4518
rect 10916 4499 10949 4507
rect 10916 4482 10924 4499
rect 10941 4482 10949 4499
rect 10916 4474 10949 4482
rect 11250 4483 11283 4491
rect 11250 4466 11258 4483
rect 11275 4466 11283 4483
rect 11250 4458 11283 4466
rect 11300 4441 11327 4510
rect 11450 4441 11477 4564
rect 11911 4809 11969 4817
rect 11911 4792 11947 4809
rect 11964 4792 11969 4809
rect 11911 4775 11969 4792
rect 11911 4758 11947 4775
rect 11964 4758 11969 4775
rect 11911 4741 11969 4758
rect 11911 4724 11947 4741
rect 11964 4724 11969 4741
rect 11911 4707 11969 4724
rect 11911 4690 11947 4707
rect 11964 4690 11969 4707
rect 11911 4673 11969 4690
rect 11911 4656 11947 4673
rect 11964 4656 11969 4673
rect 11911 4639 11969 4656
rect 11911 4622 11947 4639
rect 11964 4622 11969 4639
rect 11911 4614 11969 4622
rect 11986 4809 12013 4832
rect 12597 4832 12601 4851
rect 12620 4832 12624 4851
rect 11986 4792 11991 4809
rect 12008 4792 12013 4809
rect 11986 4775 12013 4792
rect 11986 4758 11991 4775
rect 12008 4758 12013 4775
rect 11986 4741 12013 4758
rect 11986 4724 11991 4741
rect 12008 4724 12013 4741
rect 11986 4707 12013 4724
rect 11986 4690 11991 4707
rect 12008 4690 12013 4707
rect 11986 4673 12013 4690
rect 11986 4656 11991 4673
rect 12008 4656 12013 4673
rect 11986 4639 12013 4656
rect 11986 4622 11991 4639
rect 12008 4622 12013 4639
rect 11986 4614 12013 4622
rect 12030 4809 12088 4817
rect 12030 4792 12035 4809
rect 12052 4792 12088 4809
rect 12030 4775 12088 4792
rect 12030 4758 12035 4775
rect 12052 4758 12088 4775
rect 12030 4741 12088 4758
rect 12030 4724 12035 4741
rect 12052 4724 12088 4741
rect 12030 4707 12088 4724
rect 12030 4690 12035 4707
rect 12052 4690 12088 4707
rect 12030 4673 12088 4690
rect 12030 4656 12035 4673
rect 12052 4656 12088 4673
rect 12030 4639 12088 4656
rect 12030 4622 12035 4639
rect 12052 4622 12088 4639
rect 12030 4614 12088 4622
rect 11861 4537 11894 4545
rect 11861 4520 11869 4537
rect 11886 4520 11894 4537
rect 11861 4512 11894 4520
rect 11911 4527 11938 4614
rect 11960 4589 11993 4597
rect 11960 4572 11968 4589
rect 11985 4581 11993 4589
rect 12061 4581 12088 4614
rect 11985 4572 12088 4581
rect 11960 4564 12088 4572
rect 12006 4535 12039 4543
rect 12006 4527 12014 4535
rect 11911 4518 12014 4527
rect 12031 4518 12039 4535
rect 11911 4510 12039 4518
rect 11494 4499 11527 4507
rect 11494 4482 11502 4499
rect 11519 4482 11527 4499
rect 11494 4474 11527 4482
rect 11861 4483 11894 4491
rect 11861 4466 11869 4483
rect 11886 4466 11894 4483
rect 11861 4458 11894 4466
rect 11911 4441 11938 4510
rect 12061 4441 12088 4564
rect 12522 4809 12580 4817
rect 12522 4792 12558 4809
rect 12575 4792 12580 4809
rect 12522 4775 12580 4792
rect 12522 4758 12558 4775
rect 12575 4758 12580 4775
rect 12522 4741 12580 4758
rect 12522 4724 12558 4741
rect 12575 4724 12580 4741
rect 12522 4707 12580 4724
rect 12522 4690 12558 4707
rect 12575 4690 12580 4707
rect 12522 4673 12580 4690
rect 12522 4656 12558 4673
rect 12575 4656 12580 4673
rect 12522 4639 12580 4656
rect 12522 4622 12558 4639
rect 12575 4622 12580 4639
rect 12522 4614 12580 4622
rect 12597 4809 12624 4832
rect 12597 4792 12602 4809
rect 12619 4792 12624 4809
rect 12597 4775 12624 4792
rect 12597 4758 12602 4775
rect 12619 4758 12624 4775
rect 12597 4741 12624 4758
rect 12597 4724 12602 4741
rect 12619 4724 12624 4741
rect 12597 4707 12624 4724
rect 12597 4690 12602 4707
rect 12619 4690 12624 4707
rect 12597 4673 12624 4690
rect 12597 4656 12602 4673
rect 12619 4656 12624 4673
rect 12597 4639 12624 4656
rect 12597 4622 12602 4639
rect 12619 4622 12624 4639
rect 12597 4614 12624 4622
rect 12641 4809 12699 4817
rect 12641 4792 12646 4809
rect 12663 4792 12699 4809
rect 12641 4775 12699 4792
rect 12641 4758 12646 4775
rect 12663 4758 12699 4775
rect 12641 4741 12699 4758
rect 12641 4724 12646 4741
rect 12663 4724 12699 4741
rect 12641 4707 12699 4724
rect 12641 4690 12646 4707
rect 12663 4690 12699 4707
rect 12641 4673 12699 4690
rect 12641 4656 12646 4673
rect 12663 4656 12699 4673
rect 12641 4639 12699 4656
rect 12641 4622 12646 4639
rect 12663 4622 12699 4639
rect 12641 4614 12699 4622
rect 12472 4537 12505 4545
rect 12472 4520 12480 4537
rect 12497 4520 12505 4537
rect 12472 4512 12505 4520
rect 12522 4527 12549 4614
rect 12571 4589 12604 4597
rect 12571 4572 12579 4589
rect 12596 4581 12604 4589
rect 12672 4581 12699 4614
rect 12596 4572 12699 4581
rect 12571 4564 12699 4572
rect 12617 4535 12650 4543
rect 12617 4527 12625 4535
rect 12522 4518 12625 4527
rect 12642 4518 12650 4535
rect 12522 4510 12650 4518
rect 12105 4499 12138 4507
rect 12105 4482 12113 4499
rect 12130 4482 12138 4499
rect 12105 4474 12138 4482
rect 12472 4483 12505 4491
rect 12472 4466 12480 4483
rect 12497 4466 12505 4483
rect 12472 4458 12505 4466
rect 12522 4441 12549 4510
rect 12672 4441 12699 4564
rect 12716 4499 12749 4507
rect 12716 4482 12724 4499
rect 12741 4482 12749 4499
rect 12716 4474 12749 4482
rect 9451 4433 9478 4441
rect 9451 4416 9456 4433
rect 9473 4416 9478 4433
rect 9451 4399 9478 4416
rect 9451 4382 9456 4399
rect 9473 4382 9478 4399
rect 9451 4365 9478 4382
rect 9451 4348 9456 4365
rect 9473 4348 9478 4365
rect 9451 4340 9478 4348
rect 9500 4433 9558 4441
rect 9500 4416 9536 4433
rect 9553 4416 9558 4433
rect 9500 4399 9558 4416
rect 9500 4382 9536 4399
rect 9553 4382 9558 4399
rect 9500 4365 9558 4382
rect 9500 4348 9536 4365
rect 9553 4348 9558 4365
rect 9500 4340 9558 4348
rect 9575 4433 9602 4441
rect 9575 4416 9580 4433
rect 9597 4416 9602 4433
rect 9575 4399 9602 4416
rect 9575 4382 9580 4399
rect 9597 4382 9602 4399
rect 9575 4365 9602 4382
rect 9575 4348 9580 4365
rect 9597 4348 9602 4365
rect 9575 4325 9602 4348
rect 9619 4433 9677 4441
rect 9619 4416 9624 4433
rect 9641 4416 9677 4433
rect 9619 4399 9677 4416
rect 9619 4382 9624 4399
rect 9641 4382 9677 4399
rect 9619 4365 9677 4382
rect 9619 4348 9624 4365
rect 9641 4348 9677 4365
rect 9619 4340 9677 4348
rect 9699 4433 9726 4441
rect 9699 4416 9704 4433
rect 9721 4416 9726 4433
rect 9699 4399 9726 4416
rect 9699 4382 9704 4399
rect 9721 4382 9726 4399
rect 9699 4365 9726 4382
rect 9699 4348 9704 4365
rect 9721 4348 9726 4365
rect 9699 4340 9726 4348
rect 10062 4433 10089 4441
rect 10062 4416 10067 4433
rect 10084 4416 10089 4433
rect 10062 4399 10089 4416
rect 10062 4382 10067 4399
rect 10084 4382 10089 4399
rect 10062 4365 10089 4382
rect 10062 4348 10067 4365
rect 10084 4348 10089 4365
rect 10062 4340 10089 4348
rect 10111 4433 10169 4441
rect 10111 4416 10147 4433
rect 10164 4416 10169 4433
rect 10111 4399 10169 4416
rect 10111 4382 10147 4399
rect 10164 4382 10169 4399
rect 10111 4365 10169 4382
rect 10111 4348 10147 4365
rect 10164 4348 10169 4365
rect 10111 4340 10169 4348
rect 10186 4433 10213 4441
rect 10186 4416 10191 4433
rect 10208 4416 10213 4433
rect 10186 4399 10213 4416
rect 10186 4382 10191 4399
rect 10208 4382 10213 4399
rect 10186 4365 10213 4382
rect 10186 4348 10191 4365
rect 10208 4348 10213 4365
rect 9575 4306 9579 4325
rect 9598 4306 9602 4325
rect 10186 4325 10213 4348
rect 10230 4433 10288 4441
rect 10230 4416 10235 4433
rect 10252 4416 10288 4433
rect 10230 4399 10288 4416
rect 10230 4382 10235 4399
rect 10252 4382 10288 4399
rect 10230 4365 10288 4382
rect 10230 4348 10235 4365
rect 10252 4348 10288 4365
rect 10230 4340 10288 4348
rect 10310 4433 10337 4441
rect 10310 4416 10315 4433
rect 10332 4416 10337 4433
rect 10310 4399 10337 4416
rect 10310 4382 10315 4399
rect 10332 4382 10337 4399
rect 10310 4365 10337 4382
rect 10310 4348 10315 4365
rect 10332 4348 10337 4365
rect 10310 4340 10337 4348
rect 10673 4433 10700 4441
rect 10673 4416 10678 4433
rect 10695 4416 10700 4433
rect 10673 4399 10700 4416
rect 10673 4382 10678 4399
rect 10695 4382 10700 4399
rect 10673 4365 10700 4382
rect 10673 4348 10678 4365
rect 10695 4348 10700 4365
rect 10673 4340 10700 4348
rect 10722 4433 10780 4441
rect 10722 4416 10758 4433
rect 10775 4416 10780 4433
rect 10722 4399 10780 4416
rect 10722 4382 10758 4399
rect 10775 4382 10780 4399
rect 10722 4365 10780 4382
rect 10722 4348 10758 4365
rect 10775 4348 10780 4365
rect 10722 4340 10780 4348
rect 10797 4433 10824 4441
rect 10797 4416 10802 4433
rect 10819 4416 10824 4433
rect 10797 4399 10824 4416
rect 10797 4382 10802 4399
rect 10819 4382 10824 4399
rect 10797 4365 10824 4382
rect 10797 4348 10802 4365
rect 10819 4348 10824 4365
rect 10186 4306 10190 4325
rect 10209 4306 10213 4325
rect 10797 4325 10824 4348
rect 10841 4433 10899 4441
rect 10841 4416 10846 4433
rect 10863 4416 10899 4433
rect 10841 4399 10899 4416
rect 10841 4382 10846 4399
rect 10863 4382 10899 4399
rect 10841 4365 10899 4382
rect 10841 4348 10846 4365
rect 10863 4348 10899 4365
rect 10841 4340 10899 4348
rect 10921 4433 10948 4441
rect 10921 4416 10926 4433
rect 10943 4416 10948 4433
rect 10921 4399 10948 4416
rect 10921 4382 10926 4399
rect 10943 4382 10948 4399
rect 10921 4365 10948 4382
rect 10921 4348 10926 4365
rect 10943 4348 10948 4365
rect 10921 4340 10948 4348
rect 11251 4433 11278 4441
rect 11251 4416 11256 4433
rect 11273 4416 11278 4433
rect 11251 4399 11278 4416
rect 11251 4382 11256 4399
rect 11273 4382 11278 4399
rect 11251 4365 11278 4382
rect 11251 4348 11256 4365
rect 11273 4348 11278 4365
rect 11251 4340 11278 4348
rect 11300 4433 11358 4441
rect 11300 4416 11336 4433
rect 11353 4416 11358 4433
rect 11300 4399 11358 4416
rect 11300 4382 11336 4399
rect 11353 4382 11358 4399
rect 11300 4365 11358 4382
rect 11300 4348 11336 4365
rect 11353 4348 11358 4365
rect 11300 4340 11358 4348
rect 11375 4433 11402 4441
rect 11375 4416 11380 4433
rect 11397 4416 11402 4433
rect 11375 4399 11402 4416
rect 11375 4382 11380 4399
rect 11397 4382 11402 4399
rect 11375 4365 11402 4382
rect 11375 4348 11380 4365
rect 11397 4348 11402 4365
rect 10797 4306 10801 4325
rect 10820 4306 10824 4325
rect 11375 4325 11402 4348
rect 11419 4433 11477 4441
rect 11419 4416 11424 4433
rect 11441 4416 11477 4433
rect 11419 4399 11477 4416
rect 11419 4382 11424 4399
rect 11441 4382 11477 4399
rect 11419 4365 11477 4382
rect 11419 4348 11424 4365
rect 11441 4348 11477 4365
rect 11419 4340 11477 4348
rect 11499 4433 11526 4441
rect 11499 4416 11504 4433
rect 11521 4416 11526 4433
rect 11499 4399 11526 4416
rect 11499 4382 11504 4399
rect 11521 4382 11526 4399
rect 11499 4365 11526 4382
rect 11499 4348 11504 4365
rect 11521 4348 11526 4365
rect 11499 4340 11526 4348
rect 11862 4433 11889 4441
rect 11862 4416 11867 4433
rect 11884 4416 11889 4433
rect 11862 4399 11889 4416
rect 11862 4382 11867 4399
rect 11884 4382 11889 4399
rect 11862 4365 11889 4382
rect 11862 4348 11867 4365
rect 11884 4348 11889 4365
rect 11862 4340 11889 4348
rect 11911 4433 11969 4441
rect 11911 4416 11947 4433
rect 11964 4416 11969 4433
rect 11911 4399 11969 4416
rect 11911 4382 11947 4399
rect 11964 4382 11969 4399
rect 11911 4365 11969 4382
rect 11911 4348 11947 4365
rect 11964 4348 11969 4365
rect 11911 4340 11969 4348
rect 11986 4433 12013 4441
rect 11986 4416 11991 4433
rect 12008 4416 12013 4433
rect 11986 4399 12013 4416
rect 11986 4382 11991 4399
rect 12008 4382 12013 4399
rect 11986 4365 12013 4382
rect 11986 4348 11991 4365
rect 12008 4348 12013 4365
rect 11375 4306 11379 4325
rect 11398 4306 11402 4325
rect 11986 4325 12013 4348
rect 12030 4433 12088 4441
rect 12030 4416 12035 4433
rect 12052 4416 12088 4433
rect 12030 4399 12088 4416
rect 12030 4382 12035 4399
rect 12052 4382 12088 4399
rect 12030 4365 12088 4382
rect 12030 4348 12035 4365
rect 12052 4348 12088 4365
rect 12030 4340 12088 4348
rect 12110 4433 12137 4441
rect 12110 4416 12115 4433
rect 12132 4416 12137 4433
rect 12110 4399 12137 4416
rect 12110 4382 12115 4399
rect 12132 4382 12137 4399
rect 12110 4365 12137 4382
rect 12110 4348 12115 4365
rect 12132 4348 12137 4365
rect 12110 4340 12137 4348
rect 12473 4433 12500 4441
rect 12473 4416 12478 4433
rect 12495 4416 12500 4433
rect 12473 4399 12500 4416
rect 12473 4382 12478 4399
rect 12495 4382 12500 4399
rect 12473 4365 12500 4382
rect 12473 4348 12478 4365
rect 12495 4348 12500 4365
rect 12473 4340 12500 4348
rect 12522 4433 12580 4441
rect 12522 4416 12558 4433
rect 12575 4416 12580 4433
rect 12522 4399 12580 4416
rect 12522 4382 12558 4399
rect 12575 4382 12580 4399
rect 12522 4365 12580 4382
rect 12522 4348 12558 4365
rect 12575 4348 12580 4365
rect 12522 4340 12580 4348
rect 12597 4433 12624 4441
rect 12597 4416 12602 4433
rect 12619 4416 12624 4433
rect 12597 4399 12624 4416
rect 12597 4382 12602 4399
rect 12619 4382 12624 4399
rect 12597 4365 12624 4382
rect 12597 4348 12602 4365
rect 12619 4348 12624 4365
rect 11986 4306 11990 4325
rect 12009 4306 12013 4325
rect 12597 4325 12624 4348
rect 12641 4433 12699 4441
rect 12641 4416 12646 4433
rect 12663 4416 12699 4433
rect 12641 4399 12699 4416
rect 12641 4382 12646 4399
rect 12663 4382 12699 4399
rect 12641 4365 12699 4382
rect 12641 4348 12646 4365
rect 12663 4348 12699 4365
rect 12641 4340 12699 4348
rect 12721 4433 12748 4441
rect 12721 4416 12726 4433
rect 12743 4416 12748 4433
rect 12721 4399 12748 4416
rect 12721 4382 12726 4399
rect 12743 4382 12748 4399
rect 12721 4365 12748 4382
rect 12721 4348 12726 4365
rect 12743 4348 12748 4365
rect 12721 4340 12748 4348
rect 12597 4306 12601 4325
rect 12620 4306 12624 4325
<< viali >>
rect 10190 8062 10209 8081
rect 10801 8062 10820 8081
rect 10069 7750 10086 7767
rect 10168 7802 10185 7819
rect 10214 7748 10231 7765
rect 10069 7696 10086 7713
rect 11379 8062 11398 8081
rect 10680 7750 10697 7767
rect 10779 7802 10796 7819
rect 10825 7748 10842 7765
rect 10313 7712 10330 7729
rect 10680 7696 10697 7713
rect 11990 8062 12009 8081
rect 11258 7750 11275 7767
rect 11357 7802 11374 7819
rect 11403 7748 11420 7765
rect 10924 7712 10941 7729
rect 11258 7696 11275 7713
rect 12601 8062 12620 8081
rect 11869 7750 11886 7767
rect 11968 7802 11985 7819
rect 12014 7748 12031 7765
rect 11502 7712 11519 7729
rect 11869 7696 11886 7713
rect 12480 7750 12497 7767
rect 12579 7802 12596 7819
rect 12625 7748 12642 7765
rect 12113 7712 12130 7729
rect 12480 7696 12497 7713
rect 12724 7712 12741 7729
rect 10190 7536 10209 7555
rect 10801 7536 10820 7555
rect 11379 7536 11398 7555
rect 11990 7536 12009 7555
rect 12601 7536 12620 7555
rect 9579 7412 9598 7431
rect 10190 7412 10209 7431
rect 9458 7100 9475 7117
rect 9557 7152 9574 7169
rect 9603 7098 9620 7115
rect 9458 7046 9475 7063
rect 10801 7412 10820 7431
rect 10069 7100 10086 7117
rect 10168 7152 10185 7169
rect 10214 7098 10231 7115
rect 9702 7062 9719 7079
rect 10069 7046 10086 7063
rect 11379 7412 11398 7431
rect 10680 7100 10697 7117
rect 10779 7152 10796 7169
rect 10825 7098 10842 7115
rect 10313 7062 10330 7079
rect 10680 7046 10697 7063
rect 11990 7412 12009 7431
rect 11258 7100 11275 7117
rect 11357 7152 11374 7169
rect 11403 7098 11420 7115
rect 10924 7062 10941 7079
rect 11258 7046 11275 7063
rect 12601 7412 12620 7431
rect 11869 7100 11886 7117
rect 11968 7152 11985 7169
rect 12014 7098 12031 7115
rect 11502 7062 11519 7079
rect 11869 7046 11886 7063
rect 12480 7100 12497 7117
rect 12579 7152 12596 7169
rect 12625 7098 12642 7115
rect 12113 7062 12130 7079
rect 12480 7046 12497 7063
rect 12724 7062 12741 7079
rect 9579 6886 9598 6905
rect 10190 6886 10209 6905
rect 10801 6886 10820 6905
rect 11379 6886 11398 6905
rect 11990 6886 12009 6905
rect 12601 6886 12620 6905
rect 9579 6772 9598 6791
rect 10190 6772 10209 6791
rect 9458 6460 9475 6477
rect 9557 6512 9574 6529
rect 9603 6458 9620 6475
rect 9458 6406 9475 6423
rect 10801 6772 10820 6791
rect 10069 6460 10086 6477
rect 10168 6512 10185 6529
rect 10214 6458 10231 6475
rect 9702 6422 9719 6439
rect 10069 6406 10086 6423
rect 11379 6772 11398 6791
rect 10680 6460 10697 6477
rect 10779 6512 10796 6529
rect 10825 6458 10842 6475
rect 10313 6422 10330 6439
rect 10680 6406 10697 6423
rect 11990 6772 12009 6791
rect 11258 6460 11275 6477
rect 11357 6512 11374 6529
rect 11403 6458 11420 6475
rect 10924 6422 10941 6439
rect 11258 6406 11275 6423
rect 12601 6772 12620 6791
rect 11869 6460 11886 6477
rect 11968 6512 11985 6529
rect 12014 6458 12031 6475
rect 11502 6422 11519 6439
rect 11869 6406 11886 6423
rect 12480 6460 12497 6477
rect 12579 6512 12596 6529
rect 12625 6458 12642 6475
rect 12113 6422 12130 6439
rect 12480 6406 12497 6423
rect 12724 6422 12741 6439
rect 9579 6246 9598 6265
rect 10190 6246 10209 6265
rect 10801 6246 10820 6265
rect 11379 6246 11398 6265
rect 11990 6246 12009 6265
rect 12601 6246 12620 6265
rect 9579 6122 9598 6141
rect 10190 6122 10209 6141
rect 9458 5810 9475 5827
rect 9557 5862 9574 5879
rect 9603 5808 9620 5825
rect 9458 5756 9475 5773
rect 10801 6122 10820 6141
rect 10069 5810 10086 5827
rect 10168 5862 10185 5879
rect 10214 5808 10231 5825
rect 9702 5772 9719 5789
rect 10069 5756 10086 5773
rect 11379 6122 11398 6141
rect 10680 5810 10697 5827
rect 10779 5862 10796 5879
rect 10825 5808 10842 5825
rect 10313 5772 10330 5789
rect 10680 5756 10697 5773
rect 11990 6122 12009 6141
rect 11258 5810 11275 5827
rect 11357 5862 11374 5879
rect 11403 5808 11420 5825
rect 10924 5772 10941 5789
rect 11258 5756 11275 5773
rect 12601 6122 12620 6141
rect 11869 5810 11886 5827
rect 11968 5862 11985 5879
rect 12014 5808 12031 5825
rect 11502 5772 11519 5789
rect 11869 5756 11886 5773
rect 12480 5810 12497 5827
rect 12579 5862 12596 5879
rect 12625 5808 12642 5825
rect 12113 5772 12130 5789
rect 12480 5756 12497 5773
rect 12724 5772 12741 5789
rect 9579 5596 9598 5615
rect 10190 5596 10209 5615
rect 10801 5596 10820 5615
rect 11379 5596 11398 5615
rect 11990 5596 12009 5615
rect 12601 5596 12620 5615
rect 9579 5472 9598 5491
rect 10190 5472 10209 5491
rect 9458 5160 9475 5177
rect 9557 5212 9574 5229
rect 9603 5158 9620 5175
rect 9458 5106 9475 5123
rect 10801 5472 10820 5491
rect 10069 5160 10086 5177
rect 10168 5212 10185 5229
rect 10214 5158 10231 5175
rect 9702 5122 9719 5139
rect 10069 5106 10086 5123
rect 11379 5472 11398 5491
rect 10680 5160 10697 5177
rect 10779 5212 10796 5229
rect 10825 5158 10842 5175
rect 10313 5122 10330 5139
rect 10680 5106 10697 5123
rect 11990 5472 12009 5491
rect 11258 5160 11275 5177
rect 11357 5212 11374 5229
rect 11403 5158 11420 5175
rect 10924 5122 10941 5139
rect 11258 5106 11275 5123
rect 12601 5472 12620 5491
rect 11869 5160 11886 5177
rect 11968 5212 11985 5229
rect 12014 5158 12031 5175
rect 11502 5122 11519 5139
rect 11869 5106 11886 5123
rect 12480 5160 12497 5177
rect 12579 5212 12596 5229
rect 12625 5158 12642 5175
rect 12113 5122 12130 5139
rect 12480 5106 12497 5123
rect 12724 5122 12741 5139
rect 9579 4946 9598 4965
rect 10190 4946 10209 4965
rect 10801 4946 10820 4965
rect 11379 4946 11398 4965
rect 11990 4946 12009 4965
rect 12601 4946 12620 4965
rect 9579 4832 9598 4851
rect 10190 4832 10209 4851
rect 9458 4520 9475 4537
rect 9557 4572 9574 4589
rect 9603 4518 9620 4535
rect 9458 4466 9475 4483
rect 10801 4832 10820 4851
rect 10069 4520 10086 4537
rect 10168 4572 10185 4589
rect 10214 4518 10231 4535
rect 9702 4482 9719 4499
rect 10069 4466 10086 4483
rect 11379 4832 11398 4851
rect 10680 4520 10697 4537
rect 10779 4572 10796 4589
rect 10825 4518 10842 4535
rect 10313 4482 10330 4499
rect 10680 4466 10697 4483
rect 11990 4832 12009 4851
rect 11258 4520 11275 4537
rect 11357 4572 11374 4589
rect 11403 4518 11420 4535
rect 10924 4482 10941 4499
rect 11258 4466 11275 4483
rect 12601 4832 12620 4851
rect 11869 4520 11886 4537
rect 11968 4572 11985 4589
rect 12014 4518 12031 4535
rect 11502 4482 11519 4499
rect 11869 4466 11886 4483
rect 12480 4520 12497 4537
rect 12579 4572 12596 4589
rect 12625 4518 12642 4535
rect 12113 4482 12130 4499
rect 12480 4466 12497 4483
rect 12724 4482 12741 4499
rect 9579 4306 9598 4325
rect 10190 4306 10209 4325
rect 10801 4306 10820 4325
rect 11379 4306 11398 4325
rect 11990 4306 12009 4325
rect 12601 4306 12620 4325
<< metal1 >>
rect 9280 8081 12891 8096
rect 9280 8062 10190 8081
rect 10209 8062 10801 8081
rect 10820 8062 11379 8081
rect 11398 8062 11990 8081
rect 12009 8062 12601 8081
rect 12620 8062 12891 8081
rect 9280 8047 12891 8062
rect 9518 7824 9582 7827
rect 9518 7797 9521 7824
rect 9548 7797 9582 7824
rect 9518 7794 9582 7797
rect 10160 7819 10193 7827
rect 10160 7802 10168 7819
rect 10185 7802 10193 7819
rect 10160 7794 10193 7802
rect 10771 7819 10804 7827
rect 10771 7802 10779 7819
rect 10796 7802 10804 7819
rect 10771 7794 10804 7802
rect 11318 7824 11382 7827
rect 11318 7797 11321 7824
rect 11348 7819 11382 7824
rect 11348 7802 11357 7819
rect 11374 7802 11382 7819
rect 11348 7797 11382 7802
rect 11318 7794 11382 7797
rect 11960 7819 11993 7827
rect 11960 7802 11968 7819
rect 11985 7802 11993 7819
rect 11960 7794 11993 7802
rect 12571 7819 12604 7827
rect 12571 7802 12579 7819
rect 12596 7802 12604 7819
rect 12571 7794 12604 7802
rect 9302 7771 9483 7775
rect 9302 7745 9305 7771
rect 9331 7745 9483 7771
rect 9302 7742 9483 7745
rect 9595 7770 9661 7773
rect 9595 7743 9631 7770
rect 9658 7743 9661 7770
rect 9595 7740 9661 7743
rect 9913 7771 10094 7775
rect 9913 7745 9916 7771
rect 9942 7767 10094 7771
rect 9942 7750 10069 7767
rect 10086 7750 10094 7767
rect 9942 7745 10094 7750
rect 9913 7742 10094 7745
rect 10206 7765 10239 7773
rect 10206 7748 10214 7765
rect 10231 7748 10239 7765
rect 10206 7740 10239 7748
rect 10524 7771 10705 7775
rect 10524 7745 10527 7771
rect 10553 7767 10705 7771
rect 10553 7750 10680 7767
rect 10697 7750 10705 7767
rect 10553 7745 10705 7750
rect 10524 7742 10705 7745
rect 10817 7765 10850 7773
rect 10817 7748 10825 7765
rect 10842 7748 10850 7765
rect 10817 7740 10850 7748
rect 11102 7771 11283 7775
rect 11102 7745 11105 7771
rect 11131 7767 11283 7771
rect 11131 7750 11258 7767
rect 11275 7750 11283 7767
rect 11131 7745 11283 7750
rect 11102 7742 11283 7745
rect 11395 7770 11461 7773
rect 11395 7765 11431 7770
rect 11395 7748 11403 7765
rect 11420 7748 11431 7765
rect 11395 7743 11431 7748
rect 11458 7743 11461 7770
rect 11395 7740 11461 7743
rect 11713 7771 11894 7775
rect 11713 7745 11716 7771
rect 11742 7767 11894 7771
rect 11742 7750 11869 7767
rect 11886 7750 11894 7767
rect 11742 7745 11894 7750
rect 11713 7742 11894 7745
rect 12006 7765 12039 7773
rect 12006 7748 12014 7765
rect 12031 7748 12039 7765
rect 12006 7740 12039 7748
rect 12324 7771 12505 7775
rect 12324 7745 12327 7771
rect 12353 7767 12505 7771
rect 12353 7750 12480 7767
rect 12497 7750 12505 7767
rect 12353 7745 12505 7750
rect 12324 7742 12505 7745
rect 12617 7765 12650 7773
rect 12617 7748 12625 7765
rect 12642 7748 12650 7765
rect 12617 7740 12650 7748
rect 9694 7733 9805 7737
rect 9402 7717 9483 7721
rect 9402 7691 9405 7717
rect 9431 7691 9483 7717
rect 9694 7707 9775 7733
rect 9801 7707 9805 7733
rect 10305 7733 10416 7737
rect 10305 7729 10386 7733
rect 9694 7704 9805 7707
rect 10013 7717 10094 7721
rect 9402 7688 9483 7691
rect 10013 7691 10016 7717
rect 10042 7713 10094 7717
rect 10042 7696 10069 7713
rect 10086 7696 10094 7713
rect 10305 7712 10313 7729
rect 10330 7712 10386 7729
rect 10305 7707 10386 7712
rect 10412 7707 10416 7733
rect 10916 7733 11027 7737
rect 10916 7729 10997 7733
rect 10305 7704 10416 7707
rect 10624 7717 10705 7721
rect 10042 7691 10094 7696
rect 10013 7688 10094 7691
rect 10624 7691 10627 7717
rect 10653 7713 10705 7717
rect 10653 7696 10680 7713
rect 10697 7696 10705 7713
rect 10916 7712 10924 7729
rect 10941 7712 10997 7729
rect 10916 7707 10997 7712
rect 11023 7707 11027 7733
rect 11494 7733 11605 7737
rect 11494 7729 11575 7733
rect 10916 7704 11027 7707
rect 11202 7717 11283 7721
rect 10653 7691 10705 7696
rect 10624 7688 10705 7691
rect 11202 7691 11205 7717
rect 11231 7713 11283 7717
rect 11231 7696 11258 7713
rect 11275 7696 11283 7713
rect 11494 7712 11502 7729
rect 11519 7712 11575 7729
rect 11494 7707 11575 7712
rect 11601 7707 11605 7733
rect 12105 7733 12216 7737
rect 12105 7729 12186 7733
rect 11494 7704 11605 7707
rect 11813 7717 11894 7721
rect 11231 7691 11283 7696
rect 11202 7688 11283 7691
rect 11813 7691 11816 7717
rect 11842 7713 11894 7717
rect 11842 7696 11869 7713
rect 11886 7696 11894 7713
rect 12105 7712 12113 7729
rect 12130 7712 12186 7729
rect 12105 7707 12186 7712
rect 12212 7707 12216 7733
rect 12716 7733 12827 7737
rect 12716 7729 12797 7733
rect 12105 7704 12216 7707
rect 12424 7717 12505 7721
rect 11842 7691 11894 7696
rect 11813 7688 11894 7691
rect 12424 7691 12427 7717
rect 12453 7713 12505 7717
rect 12453 7696 12480 7713
rect 12497 7696 12505 7713
rect 12716 7712 12724 7729
rect 12741 7712 12797 7729
rect 12716 7707 12797 7712
rect 12823 7707 12827 7733
rect 12716 7704 12827 7707
rect 12453 7691 12505 7696
rect 12424 7688 12505 7691
rect 9247 7555 12891 7570
rect 9247 7536 10190 7555
rect 10209 7536 10801 7555
rect 10820 7536 11379 7555
rect 11398 7536 11990 7555
rect 12009 7536 12601 7555
rect 12620 7536 12891 7555
rect 9247 7521 12891 7536
rect 9261 7431 12891 7446
rect 9261 7412 9579 7431
rect 9598 7412 10190 7431
rect 10209 7412 10801 7431
rect 10820 7412 11379 7431
rect 11398 7412 11990 7431
rect 12009 7412 12601 7431
rect 12620 7412 12891 7431
rect 9261 7397 12891 7412
rect 9516 7174 9582 7177
rect 9516 7147 9519 7174
rect 9546 7169 9582 7174
rect 9546 7152 9557 7169
rect 9574 7152 9582 7169
rect 9546 7147 9582 7152
rect 9516 7144 9582 7147
rect 10127 7173 10193 7177
rect 10127 7146 10133 7173
rect 10160 7169 10193 7173
rect 10160 7152 10168 7169
rect 10185 7152 10193 7169
rect 10160 7146 10193 7152
rect 10127 7144 10193 7146
rect 10738 7173 10804 7177
rect 10738 7146 10743 7173
rect 10770 7169 10804 7173
rect 10770 7152 10779 7169
rect 10796 7152 10804 7169
rect 10770 7146 10804 7152
rect 10738 7144 10804 7146
rect 11316 7174 11382 7177
rect 11316 7147 11319 7174
rect 11346 7169 11382 7174
rect 11346 7152 11357 7169
rect 11374 7152 11382 7169
rect 11346 7147 11382 7152
rect 11316 7144 11382 7147
rect 11927 7173 11993 7177
rect 11927 7146 11933 7173
rect 11960 7169 11993 7173
rect 11960 7152 11968 7169
rect 11985 7152 11993 7169
rect 11960 7146 11993 7152
rect 11927 7144 11993 7146
rect 12538 7173 12604 7177
rect 12538 7146 12543 7173
rect 12570 7169 12604 7173
rect 12570 7152 12579 7169
rect 12596 7152 12604 7169
rect 12570 7146 12604 7152
rect 12538 7144 12604 7146
rect 9302 7121 9483 7125
rect 9302 7095 9305 7121
rect 9331 7117 9483 7121
rect 9331 7100 9458 7117
rect 9475 7100 9483 7117
rect 9331 7095 9483 7100
rect 9302 7092 9483 7095
rect 9595 7120 9661 7123
rect 9595 7115 9631 7120
rect 9595 7098 9603 7115
rect 9620 7098 9631 7115
rect 9595 7093 9631 7098
rect 9658 7093 9661 7120
rect 9595 7090 9661 7093
rect 9913 7121 10094 7125
rect 9913 7095 9916 7121
rect 9942 7117 10094 7121
rect 9942 7100 10069 7117
rect 10086 7100 10094 7117
rect 9942 7095 10094 7100
rect 9913 7092 10094 7095
rect 10206 7120 10266 7123
rect 10206 7115 10239 7120
rect 10206 7098 10214 7115
rect 10231 7098 10239 7115
rect 10206 7093 10239 7098
rect 10206 7090 10266 7093
rect 10524 7121 10705 7125
rect 10524 7095 10527 7121
rect 10553 7117 10705 7121
rect 10553 7100 10680 7117
rect 10697 7100 10705 7117
rect 10553 7095 10705 7100
rect 10524 7092 10705 7095
rect 10817 7120 10882 7123
rect 10817 7115 10851 7120
rect 10817 7098 10825 7115
rect 10842 7098 10851 7115
rect 10817 7093 10851 7098
rect 10878 7093 10882 7120
rect 10817 7090 10882 7093
rect 11102 7121 11283 7125
rect 11102 7095 11105 7121
rect 11131 7117 11283 7121
rect 11131 7100 11258 7117
rect 11275 7100 11283 7117
rect 11131 7095 11283 7100
rect 11102 7092 11283 7095
rect 11395 7120 11461 7123
rect 11395 7115 11431 7120
rect 11395 7098 11403 7115
rect 11420 7098 11431 7115
rect 11395 7093 11431 7098
rect 11458 7093 11461 7120
rect 11395 7090 11461 7093
rect 11713 7121 11894 7125
rect 11713 7095 11716 7121
rect 11742 7117 11894 7121
rect 11742 7100 11869 7117
rect 11886 7100 11894 7117
rect 11742 7095 11894 7100
rect 11713 7092 11894 7095
rect 12006 7120 12066 7123
rect 12006 7115 12039 7120
rect 12006 7098 12014 7115
rect 12031 7098 12039 7115
rect 12006 7093 12039 7098
rect 12006 7090 12066 7093
rect 12324 7121 12505 7125
rect 12324 7095 12327 7121
rect 12353 7117 12505 7121
rect 12353 7100 12480 7117
rect 12497 7100 12505 7117
rect 12353 7095 12505 7100
rect 12324 7092 12505 7095
rect 12617 7120 12682 7123
rect 12617 7115 12651 7120
rect 12617 7098 12625 7115
rect 12642 7098 12651 7115
rect 12617 7093 12651 7098
rect 12678 7093 12682 7120
rect 12617 7090 12682 7093
rect 10234 7089 10266 7090
rect 12034 7089 12066 7090
rect 9694 7083 9805 7087
rect 9694 7079 9775 7083
rect 9402 7067 9483 7071
rect 9402 7041 9405 7067
rect 9431 7063 9483 7067
rect 9431 7046 9458 7063
rect 9475 7046 9483 7063
rect 9694 7062 9702 7079
rect 9719 7062 9775 7079
rect 9694 7057 9775 7062
rect 9801 7057 9805 7083
rect 10305 7083 10416 7087
rect 10305 7079 10386 7083
rect 9694 7054 9805 7057
rect 10013 7067 10094 7071
rect 9431 7041 9483 7046
rect 9402 7038 9483 7041
rect 10013 7041 10016 7067
rect 10042 7063 10094 7067
rect 10042 7046 10069 7063
rect 10086 7046 10094 7063
rect 10305 7062 10313 7079
rect 10330 7062 10386 7079
rect 10305 7057 10386 7062
rect 10412 7057 10416 7083
rect 10916 7083 11027 7087
rect 10916 7079 10997 7083
rect 10305 7054 10416 7057
rect 10624 7067 10705 7071
rect 10042 7041 10094 7046
rect 10013 7038 10094 7041
rect 10624 7041 10627 7067
rect 10653 7063 10705 7067
rect 10653 7046 10680 7063
rect 10697 7046 10705 7063
rect 10916 7062 10924 7079
rect 10941 7062 10997 7079
rect 10916 7057 10997 7062
rect 11023 7057 11027 7083
rect 11494 7083 11605 7087
rect 11494 7079 11575 7083
rect 10916 7054 11027 7057
rect 11202 7067 11283 7071
rect 10653 7041 10705 7046
rect 10624 7038 10705 7041
rect 11202 7041 11205 7067
rect 11231 7063 11283 7067
rect 11231 7046 11258 7063
rect 11275 7046 11283 7063
rect 11494 7062 11502 7079
rect 11519 7062 11575 7079
rect 11494 7057 11575 7062
rect 11601 7057 11605 7083
rect 12105 7083 12216 7087
rect 12105 7079 12186 7083
rect 11494 7054 11605 7057
rect 11813 7067 11894 7071
rect 11231 7041 11283 7046
rect 11202 7038 11283 7041
rect 11813 7041 11816 7067
rect 11842 7063 11894 7067
rect 11842 7046 11869 7063
rect 11886 7046 11894 7063
rect 12105 7062 12113 7079
rect 12130 7062 12186 7079
rect 12105 7057 12186 7062
rect 12212 7057 12216 7083
rect 12716 7083 12827 7087
rect 12716 7079 12797 7083
rect 12105 7054 12216 7057
rect 12424 7067 12505 7071
rect 11842 7041 11894 7046
rect 11813 7038 11894 7041
rect 12424 7041 12427 7067
rect 12453 7063 12505 7067
rect 12453 7046 12480 7063
rect 12497 7046 12505 7063
rect 12716 7062 12724 7079
rect 12741 7062 12797 7079
rect 12716 7057 12797 7062
rect 12823 7057 12827 7083
rect 12716 7054 12827 7057
rect 12453 7041 12505 7046
rect 12424 7038 12505 7041
rect 9235 6905 12891 6920
rect 9235 6886 9579 6905
rect 9598 6886 10190 6905
rect 10209 6886 10801 6905
rect 10820 6886 11379 6905
rect 11398 6886 11990 6905
rect 12009 6886 12601 6905
rect 12620 6886 12891 6905
rect 9235 6871 12891 6886
rect 9253 6791 12891 6806
rect 9253 6772 9579 6791
rect 9598 6772 10190 6791
rect 10209 6772 10801 6791
rect 10820 6772 11379 6791
rect 11398 6772 11990 6791
rect 12009 6772 12601 6791
rect 12620 6772 12891 6791
rect 9253 6757 12891 6772
rect 9516 6534 9582 6537
rect 9516 6507 9519 6534
rect 9546 6529 9582 6534
rect 9546 6512 9557 6529
rect 9574 6512 9582 6529
rect 9546 6507 9582 6512
rect 9516 6504 9582 6507
rect 10128 6534 10193 6537
rect 10128 6507 10133 6534
rect 10160 6529 10193 6534
rect 10160 6512 10168 6529
rect 10185 6512 10193 6529
rect 10160 6507 10193 6512
rect 10128 6504 10193 6507
rect 10739 6534 10804 6537
rect 10739 6507 10744 6534
rect 10771 6529 10804 6534
rect 10771 6512 10779 6529
rect 10796 6512 10804 6529
rect 10771 6507 10804 6512
rect 10739 6504 10804 6507
rect 11316 6534 11382 6537
rect 11316 6507 11319 6534
rect 11346 6529 11382 6534
rect 11346 6512 11357 6529
rect 11374 6512 11382 6529
rect 11346 6507 11382 6512
rect 11316 6504 11382 6507
rect 11928 6534 11993 6537
rect 11928 6507 11933 6534
rect 11960 6529 11993 6534
rect 11960 6512 11968 6529
rect 11985 6512 11993 6529
rect 11960 6507 11993 6512
rect 11928 6504 11993 6507
rect 12539 6534 12604 6537
rect 12539 6507 12544 6534
rect 12571 6529 12604 6534
rect 12571 6512 12579 6529
rect 12596 6512 12604 6529
rect 12571 6507 12604 6512
rect 12539 6504 12604 6507
rect 9302 6481 9483 6485
rect 9302 6455 9305 6481
rect 9331 6477 9483 6481
rect 9331 6460 9458 6477
rect 9475 6460 9483 6477
rect 9331 6455 9483 6460
rect 9302 6452 9483 6455
rect 9595 6480 9661 6483
rect 9595 6475 9631 6480
rect 9595 6458 9603 6475
rect 9620 6458 9631 6475
rect 9595 6453 9631 6458
rect 9658 6453 9661 6480
rect 9595 6450 9661 6453
rect 9913 6481 10094 6485
rect 9913 6455 9916 6481
rect 9942 6477 10094 6481
rect 9942 6460 10069 6477
rect 10086 6460 10094 6477
rect 9942 6455 10094 6460
rect 9913 6452 10094 6455
rect 10206 6480 10271 6483
rect 10206 6475 10239 6480
rect 10206 6458 10214 6475
rect 10231 6458 10239 6475
rect 10206 6453 10239 6458
rect 10266 6453 10271 6480
rect 10206 6450 10271 6453
rect 10524 6481 10705 6485
rect 10524 6455 10527 6481
rect 10553 6477 10705 6481
rect 10553 6460 10680 6477
rect 10697 6460 10705 6477
rect 10553 6455 10705 6460
rect 10524 6452 10705 6455
rect 10817 6480 10882 6483
rect 10817 6475 10850 6480
rect 10817 6458 10825 6475
rect 10842 6458 10850 6475
rect 10817 6453 10850 6458
rect 10877 6453 10882 6480
rect 10817 6450 10882 6453
rect 11102 6481 11283 6485
rect 11102 6455 11105 6481
rect 11131 6477 11283 6481
rect 11131 6460 11258 6477
rect 11275 6460 11283 6477
rect 11131 6455 11283 6460
rect 11102 6452 11283 6455
rect 11395 6480 11461 6483
rect 11395 6475 11431 6480
rect 11395 6458 11403 6475
rect 11420 6458 11431 6475
rect 11395 6453 11431 6458
rect 11458 6453 11461 6480
rect 11395 6450 11461 6453
rect 11713 6481 11894 6485
rect 11713 6455 11716 6481
rect 11742 6477 11894 6481
rect 11742 6460 11869 6477
rect 11886 6460 11894 6477
rect 11742 6455 11894 6460
rect 11713 6452 11894 6455
rect 12006 6480 12071 6483
rect 12006 6475 12039 6480
rect 12006 6458 12014 6475
rect 12031 6458 12039 6475
rect 12006 6453 12039 6458
rect 12066 6453 12071 6480
rect 12006 6450 12071 6453
rect 12324 6481 12505 6485
rect 12324 6455 12327 6481
rect 12353 6477 12505 6481
rect 12353 6460 12480 6477
rect 12497 6460 12505 6477
rect 12353 6455 12505 6460
rect 12324 6452 12505 6455
rect 12617 6480 12682 6483
rect 12617 6475 12650 6480
rect 12617 6458 12625 6475
rect 12642 6458 12650 6475
rect 12617 6453 12650 6458
rect 12677 6453 12682 6480
rect 12617 6450 12682 6453
rect 9694 6443 9805 6447
rect 9694 6439 9775 6443
rect 9402 6427 9483 6431
rect 9402 6401 9405 6427
rect 9431 6423 9483 6427
rect 9431 6406 9458 6423
rect 9475 6406 9483 6423
rect 9694 6422 9702 6439
rect 9719 6422 9775 6439
rect 9694 6417 9775 6422
rect 9801 6417 9805 6443
rect 10305 6443 10416 6447
rect 10305 6439 10386 6443
rect 9694 6414 9805 6417
rect 10013 6427 10094 6431
rect 9431 6401 9483 6406
rect 9402 6398 9483 6401
rect 10013 6401 10016 6427
rect 10042 6423 10094 6427
rect 10042 6406 10069 6423
rect 10086 6406 10094 6423
rect 10305 6422 10313 6439
rect 10330 6422 10386 6439
rect 10305 6417 10386 6422
rect 10412 6417 10416 6443
rect 10916 6443 11027 6447
rect 10916 6439 10997 6443
rect 10305 6414 10416 6417
rect 10624 6427 10705 6431
rect 10042 6401 10094 6406
rect 10013 6398 10094 6401
rect 10624 6401 10627 6427
rect 10653 6423 10705 6427
rect 10653 6406 10680 6423
rect 10697 6406 10705 6423
rect 10916 6422 10924 6439
rect 10941 6422 10997 6439
rect 10916 6417 10997 6422
rect 11023 6417 11027 6443
rect 11494 6443 11605 6447
rect 11494 6439 11575 6443
rect 10916 6414 11027 6417
rect 11202 6427 11283 6431
rect 10653 6401 10705 6406
rect 10624 6398 10705 6401
rect 11202 6401 11205 6427
rect 11231 6423 11283 6427
rect 11231 6406 11258 6423
rect 11275 6406 11283 6423
rect 11494 6422 11502 6439
rect 11519 6422 11575 6439
rect 11494 6417 11575 6422
rect 11601 6417 11605 6443
rect 12105 6443 12216 6447
rect 12105 6439 12186 6443
rect 11494 6414 11605 6417
rect 11813 6427 11894 6431
rect 11231 6401 11283 6406
rect 11202 6398 11283 6401
rect 11813 6401 11816 6427
rect 11842 6423 11894 6427
rect 11842 6406 11869 6423
rect 11886 6406 11894 6423
rect 12105 6422 12113 6439
rect 12130 6422 12186 6439
rect 12105 6417 12186 6422
rect 12212 6417 12216 6443
rect 12716 6443 12827 6447
rect 12716 6439 12797 6443
rect 12105 6414 12216 6417
rect 12424 6427 12505 6431
rect 11842 6401 11894 6406
rect 11813 6398 11894 6401
rect 12424 6401 12427 6427
rect 12453 6423 12505 6427
rect 12453 6406 12480 6423
rect 12497 6406 12505 6423
rect 12716 6422 12724 6439
rect 12741 6422 12797 6439
rect 12716 6417 12797 6422
rect 12823 6417 12827 6443
rect 12716 6414 12827 6417
rect 12453 6401 12505 6406
rect 12424 6398 12505 6401
rect 9275 6265 12891 6280
rect 9275 6246 9579 6265
rect 9598 6246 10190 6265
rect 10209 6246 10801 6265
rect 10820 6246 11379 6265
rect 11398 6246 11990 6265
rect 12009 6246 12601 6265
rect 12620 6246 12891 6265
rect 9275 6231 12891 6246
rect 9280 6141 12891 6156
rect 9280 6122 9579 6141
rect 9598 6122 10190 6141
rect 10209 6122 10801 6141
rect 10820 6122 11379 6141
rect 11398 6122 11990 6141
rect 12009 6122 12601 6141
rect 12620 6122 12891 6141
rect 9280 6107 12891 6122
rect 9518 5884 9582 5887
rect 9518 5857 9521 5884
rect 9548 5879 9582 5884
rect 9548 5862 9557 5879
rect 9574 5862 9582 5879
rect 9548 5857 9582 5862
rect 9518 5854 9582 5857
rect 10160 5879 10193 5887
rect 10160 5862 10168 5879
rect 10185 5862 10193 5879
rect 10160 5854 10193 5862
rect 10771 5879 10804 5887
rect 10771 5862 10779 5879
rect 10796 5862 10804 5879
rect 10771 5854 10804 5862
rect 11318 5884 11382 5887
rect 11318 5857 11321 5884
rect 11348 5879 11382 5884
rect 11348 5862 11357 5879
rect 11374 5862 11382 5879
rect 11348 5857 11382 5862
rect 11318 5854 11382 5857
rect 11960 5879 11993 5887
rect 11960 5862 11968 5879
rect 11985 5862 11993 5879
rect 11960 5854 11993 5862
rect 12571 5879 12604 5887
rect 12571 5862 12579 5879
rect 12596 5862 12604 5879
rect 12571 5854 12604 5862
rect 9302 5831 9483 5835
rect 9302 5805 9305 5831
rect 9331 5827 9483 5831
rect 9331 5810 9458 5827
rect 9475 5810 9483 5827
rect 9331 5805 9483 5810
rect 9302 5802 9483 5805
rect 9595 5830 9661 5833
rect 9595 5825 9631 5830
rect 9595 5808 9603 5825
rect 9620 5808 9631 5825
rect 9595 5803 9631 5808
rect 9658 5803 9661 5830
rect 9595 5800 9661 5803
rect 9913 5831 10094 5835
rect 9913 5805 9916 5831
rect 9942 5827 10094 5831
rect 9942 5810 10069 5827
rect 10086 5810 10094 5827
rect 9942 5805 10094 5810
rect 9913 5802 10094 5805
rect 10206 5825 10239 5833
rect 10206 5808 10214 5825
rect 10231 5808 10239 5825
rect 10206 5800 10239 5808
rect 10524 5831 10705 5835
rect 10524 5805 10527 5831
rect 10553 5827 10705 5831
rect 10553 5810 10680 5827
rect 10697 5810 10705 5827
rect 10553 5805 10705 5810
rect 10524 5802 10705 5805
rect 10817 5825 10850 5833
rect 10817 5808 10825 5825
rect 10842 5808 10850 5825
rect 10817 5800 10850 5808
rect 11102 5831 11283 5835
rect 11102 5805 11105 5831
rect 11131 5827 11283 5831
rect 11131 5810 11258 5827
rect 11275 5810 11283 5827
rect 11131 5805 11283 5810
rect 11102 5802 11283 5805
rect 11395 5830 11461 5833
rect 11395 5825 11431 5830
rect 11395 5808 11403 5825
rect 11420 5808 11431 5825
rect 11395 5803 11431 5808
rect 11458 5803 11461 5830
rect 11395 5800 11461 5803
rect 11713 5831 11894 5835
rect 11713 5805 11716 5831
rect 11742 5827 11894 5831
rect 11742 5810 11869 5827
rect 11886 5810 11894 5827
rect 11742 5805 11894 5810
rect 11713 5802 11894 5805
rect 12006 5825 12039 5833
rect 12006 5808 12014 5825
rect 12031 5808 12039 5825
rect 12006 5800 12039 5808
rect 12324 5831 12505 5835
rect 12324 5805 12327 5831
rect 12353 5827 12505 5831
rect 12353 5810 12480 5827
rect 12497 5810 12505 5827
rect 12353 5805 12505 5810
rect 12324 5802 12505 5805
rect 12617 5825 12650 5833
rect 12617 5808 12625 5825
rect 12642 5808 12650 5825
rect 12617 5800 12650 5808
rect 9694 5793 9805 5797
rect 9694 5789 9775 5793
rect 9402 5777 9483 5781
rect 9402 5751 9405 5777
rect 9431 5773 9483 5777
rect 9431 5756 9458 5773
rect 9475 5756 9483 5773
rect 9694 5772 9702 5789
rect 9719 5772 9775 5789
rect 9694 5767 9775 5772
rect 9801 5767 9805 5793
rect 10305 5793 10416 5797
rect 10305 5789 10386 5793
rect 9694 5764 9805 5767
rect 10013 5777 10094 5781
rect 9431 5751 9483 5756
rect 9402 5748 9483 5751
rect 10013 5751 10016 5777
rect 10042 5773 10094 5777
rect 10042 5756 10069 5773
rect 10086 5756 10094 5773
rect 10305 5772 10313 5789
rect 10330 5772 10386 5789
rect 10305 5767 10386 5772
rect 10412 5767 10416 5793
rect 10916 5793 11027 5797
rect 10916 5789 10997 5793
rect 10305 5764 10416 5767
rect 10624 5777 10705 5781
rect 10042 5751 10094 5756
rect 10013 5748 10094 5751
rect 10624 5751 10627 5777
rect 10653 5773 10705 5777
rect 10653 5756 10680 5773
rect 10697 5756 10705 5773
rect 10916 5772 10924 5789
rect 10941 5772 10997 5789
rect 10916 5767 10997 5772
rect 11023 5767 11027 5793
rect 11494 5793 11605 5797
rect 11494 5789 11575 5793
rect 10916 5764 11027 5767
rect 11202 5777 11283 5781
rect 10653 5751 10705 5756
rect 10624 5748 10705 5751
rect 11202 5751 11205 5777
rect 11231 5773 11283 5777
rect 11231 5756 11258 5773
rect 11275 5756 11283 5773
rect 11494 5772 11502 5789
rect 11519 5772 11575 5789
rect 11494 5767 11575 5772
rect 11601 5767 11605 5793
rect 12105 5793 12216 5797
rect 12105 5789 12186 5793
rect 11494 5764 11605 5767
rect 11813 5777 11894 5781
rect 11231 5751 11283 5756
rect 11202 5748 11283 5751
rect 11813 5751 11816 5777
rect 11842 5773 11894 5777
rect 11842 5756 11869 5773
rect 11886 5756 11894 5773
rect 12105 5772 12113 5789
rect 12130 5772 12186 5789
rect 12105 5767 12186 5772
rect 12212 5767 12216 5793
rect 12716 5793 12827 5797
rect 12716 5789 12797 5793
rect 12105 5764 12216 5767
rect 12424 5777 12505 5781
rect 11842 5751 11894 5756
rect 11813 5748 11894 5751
rect 12424 5751 12427 5777
rect 12453 5773 12505 5777
rect 12453 5756 12480 5773
rect 12497 5756 12505 5773
rect 12716 5772 12724 5789
rect 12741 5772 12797 5789
rect 12716 5767 12797 5772
rect 12823 5767 12827 5793
rect 12716 5764 12827 5767
rect 12453 5751 12505 5756
rect 12424 5748 12505 5751
rect 9247 5615 12891 5630
rect 9247 5596 9579 5615
rect 9598 5596 10190 5615
rect 10209 5596 10801 5615
rect 10820 5596 11379 5615
rect 11398 5596 11990 5615
rect 12009 5596 12601 5615
rect 12620 5596 12891 5615
rect 9247 5581 12891 5596
rect 9261 5491 12891 5506
rect 9261 5472 9579 5491
rect 9598 5472 10190 5491
rect 10209 5472 10801 5491
rect 10820 5472 11379 5491
rect 11398 5472 11990 5491
rect 12009 5472 12601 5491
rect 12620 5472 12891 5491
rect 9261 5457 12891 5472
rect 9516 5234 9582 5237
rect 9516 5207 9519 5234
rect 9546 5229 9582 5234
rect 9546 5212 9557 5229
rect 9574 5212 9582 5229
rect 9546 5207 9582 5212
rect 9516 5204 9582 5207
rect 10127 5233 10193 5237
rect 10127 5206 10133 5233
rect 10160 5229 10193 5233
rect 10160 5212 10168 5229
rect 10185 5212 10193 5229
rect 10160 5206 10193 5212
rect 10127 5204 10193 5206
rect 10738 5233 10804 5237
rect 10738 5206 10743 5233
rect 10770 5229 10804 5233
rect 10770 5212 10779 5229
rect 10796 5212 10804 5229
rect 10770 5206 10804 5212
rect 10738 5204 10804 5206
rect 11316 5234 11382 5237
rect 11316 5207 11319 5234
rect 11346 5229 11382 5234
rect 11346 5212 11357 5229
rect 11374 5212 11382 5229
rect 11346 5207 11382 5212
rect 11316 5204 11382 5207
rect 11927 5233 11993 5237
rect 11927 5206 11933 5233
rect 11960 5229 11993 5233
rect 11960 5212 11968 5229
rect 11985 5212 11993 5229
rect 11960 5206 11993 5212
rect 11927 5204 11993 5206
rect 12538 5233 12604 5237
rect 12538 5206 12543 5233
rect 12570 5229 12604 5233
rect 12570 5212 12579 5229
rect 12596 5212 12604 5229
rect 12570 5206 12604 5212
rect 12538 5204 12604 5206
rect 9302 5181 9483 5185
rect 9302 5155 9305 5181
rect 9331 5177 9483 5181
rect 9331 5160 9458 5177
rect 9475 5160 9483 5177
rect 9331 5155 9483 5160
rect 9302 5152 9483 5155
rect 9595 5180 9661 5183
rect 9595 5175 9631 5180
rect 9595 5158 9603 5175
rect 9620 5158 9631 5175
rect 9595 5153 9631 5158
rect 9658 5153 9661 5180
rect 9595 5150 9661 5153
rect 9913 5181 10094 5185
rect 9913 5155 9916 5181
rect 9942 5177 10094 5181
rect 9942 5160 10069 5177
rect 10086 5160 10094 5177
rect 9942 5155 10094 5160
rect 9913 5152 10094 5155
rect 10206 5180 10266 5183
rect 10206 5175 10239 5180
rect 10206 5158 10214 5175
rect 10231 5158 10239 5175
rect 10206 5153 10239 5158
rect 10206 5150 10266 5153
rect 10524 5181 10705 5185
rect 10524 5155 10527 5181
rect 10553 5177 10705 5181
rect 10553 5160 10680 5177
rect 10697 5160 10705 5177
rect 10553 5155 10705 5160
rect 10524 5152 10705 5155
rect 10817 5180 10882 5183
rect 10817 5175 10851 5180
rect 10817 5158 10825 5175
rect 10842 5158 10851 5175
rect 10817 5153 10851 5158
rect 10878 5153 10882 5180
rect 10817 5150 10882 5153
rect 11102 5181 11283 5185
rect 11102 5155 11105 5181
rect 11131 5177 11283 5181
rect 11131 5160 11258 5177
rect 11275 5160 11283 5177
rect 11131 5155 11283 5160
rect 11102 5152 11283 5155
rect 11395 5180 11461 5183
rect 11395 5175 11431 5180
rect 11395 5158 11403 5175
rect 11420 5158 11431 5175
rect 11395 5153 11431 5158
rect 11458 5153 11461 5180
rect 11395 5150 11461 5153
rect 11713 5181 11894 5185
rect 11713 5155 11716 5181
rect 11742 5177 11894 5181
rect 11742 5160 11869 5177
rect 11886 5160 11894 5177
rect 11742 5155 11894 5160
rect 11713 5152 11894 5155
rect 12006 5180 12066 5183
rect 12006 5175 12039 5180
rect 12006 5158 12014 5175
rect 12031 5158 12039 5175
rect 12006 5153 12039 5158
rect 12006 5150 12066 5153
rect 12324 5181 12505 5185
rect 12324 5155 12327 5181
rect 12353 5177 12505 5181
rect 12353 5160 12480 5177
rect 12497 5160 12505 5177
rect 12353 5155 12505 5160
rect 12324 5152 12505 5155
rect 12617 5180 12682 5183
rect 12617 5175 12651 5180
rect 12617 5158 12625 5175
rect 12642 5158 12651 5175
rect 12617 5153 12651 5158
rect 12678 5153 12682 5180
rect 12617 5150 12682 5153
rect 10234 5149 10266 5150
rect 12034 5149 12066 5150
rect 9694 5143 9805 5147
rect 9694 5139 9775 5143
rect 9402 5127 9483 5131
rect 9402 5101 9405 5127
rect 9431 5123 9483 5127
rect 9431 5106 9458 5123
rect 9475 5106 9483 5123
rect 9694 5122 9702 5139
rect 9719 5122 9775 5139
rect 9694 5117 9775 5122
rect 9801 5117 9805 5143
rect 10305 5143 10416 5147
rect 10305 5139 10386 5143
rect 9694 5114 9805 5117
rect 10013 5127 10094 5131
rect 9431 5101 9483 5106
rect 9402 5098 9483 5101
rect 10013 5101 10016 5127
rect 10042 5123 10094 5127
rect 10042 5106 10069 5123
rect 10086 5106 10094 5123
rect 10305 5122 10313 5139
rect 10330 5122 10386 5139
rect 10305 5117 10386 5122
rect 10412 5117 10416 5143
rect 10916 5143 11027 5147
rect 10916 5139 10997 5143
rect 10305 5114 10416 5117
rect 10624 5127 10705 5131
rect 10042 5101 10094 5106
rect 10013 5098 10094 5101
rect 10624 5101 10627 5127
rect 10653 5123 10705 5127
rect 10653 5106 10680 5123
rect 10697 5106 10705 5123
rect 10916 5122 10924 5139
rect 10941 5122 10997 5139
rect 10916 5117 10997 5122
rect 11023 5117 11027 5143
rect 11494 5143 11605 5147
rect 11494 5139 11575 5143
rect 10916 5114 11027 5117
rect 11202 5127 11283 5131
rect 10653 5101 10705 5106
rect 10624 5098 10705 5101
rect 11202 5101 11205 5127
rect 11231 5123 11283 5127
rect 11231 5106 11258 5123
rect 11275 5106 11283 5123
rect 11494 5122 11502 5139
rect 11519 5122 11575 5139
rect 11494 5117 11575 5122
rect 11601 5117 11605 5143
rect 12105 5143 12216 5147
rect 12105 5139 12186 5143
rect 11494 5114 11605 5117
rect 11813 5127 11894 5131
rect 11231 5101 11283 5106
rect 11202 5098 11283 5101
rect 11813 5101 11816 5127
rect 11842 5123 11894 5127
rect 11842 5106 11869 5123
rect 11886 5106 11894 5123
rect 12105 5122 12113 5139
rect 12130 5122 12186 5139
rect 12105 5117 12186 5122
rect 12212 5117 12216 5143
rect 12716 5143 12827 5147
rect 12716 5139 12797 5143
rect 12105 5114 12216 5117
rect 12424 5127 12505 5131
rect 11842 5101 11894 5106
rect 11813 5098 11894 5101
rect 12424 5101 12427 5127
rect 12453 5123 12505 5127
rect 12453 5106 12480 5123
rect 12497 5106 12505 5123
rect 12716 5122 12724 5139
rect 12741 5122 12797 5139
rect 12716 5117 12797 5122
rect 12823 5117 12827 5143
rect 12716 5114 12827 5117
rect 12453 5101 12505 5106
rect 12424 5098 12505 5101
rect 9235 4965 12891 4980
rect 9235 4946 9579 4965
rect 9598 4946 10190 4965
rect 10209 4946 10801 4965
rect 10820 4946 11379 4965
rect 11398 4946 11990 4965
rect 12009 4946 12601 4965
rect 12620 4946 12891 4965
rect 9235 4931 12891 4946
rect 9253 4851 12891 4866
rect 9253 4832 9579 4851
rect 9598 4832 10190 4851
rect 10209 4832 10801 4851
rect 10820 4832 11379 4851
rect 11398 4832 11990 4851
rect 12009 4832 12601 4851
rect 12620 4832 12891 4851
rect 9253 4817 12891 4832
rect 9516 4594 9582 4597
rect 9516 4567 9519 4594
rect 9546 4589 9582 4594
rect 9546 4572 9557 4589
rect 9574 4572 9582 4589
rect 9546 4567 9582 4572
rect 9516 4564 9582 4567
rect 10128 4594 10193 4597
rect 10128 4567 10133 4594
rect 10160 4589 10193 4594
rect 10160 4572 10168 4589
rect 10185 4572 10193 4589
rect 10160 4567 10193 4572
rect 10128 4564 10193 4567
rect 10739 4594 10804 4597
rect 10739 4567 10744 4594
rect 10771 4589 10804 4594
rect 10771 4572 10779 4589
rect 10796 4572 10804 4589
rect 10771 4567 10804 4572
rect 10739 4564 10804 4567
rect 11316 4594 11382 4597
rect 11316 4567 11319 4594
rect 11346 4589 11382 4594
rect 11346 4572 11357 4589
rect 11374 4572 11382 4589
rect 11346 4567 11382 4572
rect 11316 4564 11382 4567
rect 11928 4594 11993 4597
rect 11928 4567 11933 4594
rect 11960 4589 11993 4594
rect 11960 4572 11968 4589
rect 11985 4572 11993 4589
rect 11960 4567 11993 4572
rect 11928 4564 11993 4567
rect 12539 4594 12604 4597
rect 12539 4567 12544 4594
rect 12571 4589 12604 4594
rect 12571 4572 12579 4589
rect 12596 4572 12604 4589
rect 12571 4567 12604 4572
rect 12539 4564 12604 4567
rect 9302 4541 9483 4545
rect 9302 4515 9305 4541
rect 9331 4537 9483 4541
rect 9331 4520 9458 4537
rect 9475 4520 9483 4537
rect 9331 4515 9483 4520
rect 9302 4512 9483 4515
rect 9595 4540 9661 4543
rect 9595 4535 9631 4540
rect 9595 4518 9603 4535
rect 9620 4518 9631 4535
rect 9595 4513 9631 4518
rect 9658 4513 9661 4540
rect 9595 4510 9661 4513
rect 9913 4541 10094 4545
rect 9913 4515 9916 4541
rect 9942 4537 10094 4541
rect 9942 4520 10069 4537
rect 10086 4520 10094 4537
rect 9942 4515 10094 4520
rect 9913 4512 10094 4515
rect 10206 4540 10271 4543
rect 10206 4535 10239 4540
rect 10206 4518 10214 4535
rect 10231 4518 10239 4535
rect 10206 4513 10239 4518
rect 10266 4513 10271 4540
rect 10206 4510 10271 4513
rect 10524 4541 10705 4545
rect 10524 4515 10527 4541
rect 10553 4537 10705 4541
rect 10553 4520 10680 4537
rect 10697 4520 10705 4537
rect 10553 4515 10705 4520
rect 10524 4512 10705 4515
rect 10817 4540 10882 4543
rect 10817 4535 10850 4540
rect 10817 4518 10825 4535
rect 10842 4518 10850 4535
rect 10817 4513 10850 4518
rect 10877 4513 10882 4540
rect 10817 4510 10882 4513
rect 11102 4541 11283 4545
rect 11102 4515 11105 4541
rect 11131 4537 11283 4541
rect 11131 4520 11258 4537
rect 11275 4520 11283 4537
rect 11131 4515 11283 4520
rect 11102 4512 11283 4515
rect 11395 4540 11461 4543
rect 11395 4535 11431 4540
rect 11395 4518 11403 4535
rect 11420 4518 11431 4535
rect 11395 4513 11431 4518
rect 11458 4513 11461 4540
rect 11395 4510 11461 4513
rect 11713 4541 11894 4545
rect 11713 4515 11716 4541
rect 11742 4537 11894 4541
rect 11742 4520 11869 4537
rect 11886 4520 11894 4537
rect 11742 4515 11894 4520
rect 11713 4512 11894 4515
rect 12006 4540 12071 4543
rect 12006 4535 12039 4540
rect 12006 4518 12014 4535
rect 12031 4518 12039 4535
rect 12006 4513 12039 4518
rect 12066 4513 12071 4540
rect 12006 4510 12071 4513
rect 12324 4541 12505 4545
rect 12324 4515 12327 4541
rect 12353 4537 12505 4541
rect 12353 4520 12480 4537
rect 12497 4520 12505 4537
rect 12353 4515 12505 4520
rect 12324 4512 12505 4515
rect 12617 4540 12682 4543
rect 12617 4535 12650 4540
rect 12617 4518 12625 4535
rect 12642 4518 12650 4535
rect 12617 4513 12650 4518
rect 12677 4513 12682 4540
rect 12617 4510 12682 4513
rect 9694 4503 9805 4507
rect 9694 4499 9775 4503
rect 9402 4487 9483 4491
rect 9402 4461 9405 4487
rect 9431 4483 9483 4487
rect 9431 4466 9458 4483
rect 9475 4466 9483 4483
rect 9694 4482 9702 4499
rect 9719 4482 9775 4499
rect 9694 4477 9775 4482
rect 9801 4477 9805 4503
rect 10305 4503 10416 4507
rect 10305 4499 10386 4503
rect 9694 4474 9805 4477
rect 10013 4487 10094 4491
rect 9431 4461 9483 4466
rect 9402 4458 9483 4461
rect 10013 4461 10016 4487
rect 10042 4483 10094 4487
rect 10042 4466 10069 4483
rect 10086 4466 10094 4483
rect 10305 4482 10313 4499
rect 10330 4482 10386 4499
rect 10305 4477 10386 4482
rect 10412 4477 10416 4503
rect 10916 4503 11027 4507
rect 10916 4499 10997 4503
rect 10305 4474 10416 4477
rect 10624 4487 10705 4491
rect 10042 4461 10094 4466
rect 10013 4458 10094 4461
rect 10624 4461 10627 4487
rect 10653 4483 10705 4487
rect 10653 4466 10680 4483
rect 10697 4466 10705 4483
rect 10916 4482 10924 4499
rect 10941 4482 10997 4499
rect 10916 4477 10997 4482
rect 11023 4477 11027 4503
rect 11494 4503 11605 4507
rect 11494 4499 11575 4503
rect 10916 4474 11027 4477
rect 11202 4487 11283 4491
rect 10653 4461 10705 4466
rect 10624 4458 10705 4461
rect 11202 4461 11205 4487
rect 11231 4483 11283 4487
rect 11231 4466 11258 4483
rect 11275 4466 11283 4483
rect 11494 4482 11502 4499
rect 11519 4482 11575 4499
rect 11494 4477 11575 4482
rect 11601 4477 11605 4503
rect 12105 4503 12216 4507
rect 12105 4499 12186 4503
rect 11494 4474 11605 4477
rect 11813 4487 11894 4491
rect 11231 4461 11283 4466
rect 11202 4458 11283 4461
rect 11813 4461 11816 4487
rect 11842 4483 11894 4487
rect 11842 4466 11869 4483
rect 11886 4466 11894 4483
rect 12105 4482 12113 4499
rect 12130 4482 12186 4499
rect 12105 4477 12186 4482
rect 12212 4477 12216 4503
rect 12716 4503 12827 4507
rect 12716 4499 12797 4503
rect 12105 4474 12216 4477
rect 12424 4487 12505 4491
rect 11842 4461 11894 4466
rect 11813 4458 11894 4461
rect 12424 4461 12427 4487
rect 12453 4483 12505 4487
rect 12453 4466 12480 4483
rect 12497 4466 12505 4483
rect 12716 4482 12724 4499
rect 12741 4482 12797 4499
rect 12716 4477 12797 4482
rect 12823 4477 12827 4503
rect 12716 4474 12827 4477
rect 12453 4461 12505 4466
rect 12424 4458 12505 4461
rect 9275 4325 12891 4340
rect 9275 4306 9579 4325
rect 9598 4306 10190 4325
rect 10209 4306 10801 4325
rect 10820 4306 11379 4325
rect 11398 4306 11990 4325
rect 12009 4306 12601 4325
rect 12620 4306 12891 4325
rect 9275 4291 12891 4306
rect 975 1218 14336 1266
rect 975 1156 1025 1218
rect 600 1155 1025 1156
rect 251 1154 1025 1155
rect 100 1145 1025 1154
rect 100 1113 154 1145
rect 186 1113 1025 1145
rect 100 1105 1025 1113
rect 100 1104 400 1105
rect 13249 890 14137 915
rect 13249 850 13274 890
rect 13314 850 14137 890
rect 13249 825 14137 850
rect 14267 890 15271 915
rect 14267 850 15206 890
rect 15246 850 15271 890
rect 14267 825 15271 850
rect 400 633 14335 683
<< via1 >>
rect 9521 7797 9548 7824
rect 11321 7797 11348 7824
rect 9305 7745 9331 7771
rect 9631 7743 9658 7770
rect 9916 7745 9942 7771
rect 10527 7745 10553 7771
rect 11105 7745 11131 7771
rect 11431 7743 11458 7770
rect 11716 7745 11742 7771
rect 12327 7745 12353 7771
rect 9405 7691 9431 7717
rect 9775 7707 9801 7733
rect 10016 7691 10042 7717
rect 10386 7707 10412 7733
rect 10627 7691 10653 7717
rect 10997 7707 11023 7733
rect 11205 7691 11231 7717
rect 11575 7707 11601 7733
rect 11816 7691 11842 7717
rect 12186 7707 12212 7733
rect 12427 7691 12453 7717
rect 12797 7707 12823 7733
rect 9519 7147 9546 7174
rect 10133 7146 10160 7173
rect 10743 7146 10770 7173
rect 11319 7147 11346 7174
rect 11933 7146 11960 7173
rect 12543 7146 12570 7173
rect 9305 7095 9331 7121
rect 9631 7093 9658 7120
rect 9916 7095 9942 7121
rect 10239 7093 10266 7120
rect 10527 7095 10553 7121
rect 10851 7093 10878 7120
rect 11105 7095 11131 7121
rect 11431 7093 11458 7120
rect 11716 7095 11742 7121
rect 12039 7093 12066 7120
rect 12327 7095 12353 7121
rect 12651 7093 12678 7120
rect 9405 7041 9431 7067
rect 9775 7057 9801 7083
rect 10016 7041 10042 7067
rect 10386 7057 10412 7083
rect 10627 7041 10653 7067
rect 10997 7057 11023 7083
rect 11205 7041 11231 7067
rect 11575 7057 11601 7083
rect 11816 7041 11842 7067
rect 12186 7057 12212 7083
rect 12427 7041 12453 7067
rect 12797 7057 12823 7083
rect 9519 6507 9546 6534
rect 10133 6507 10160 6534
rect 10744 6507 10771 6534
rect 11319 6507 11346 6534
rect 11933 6507 11960 6534
rect 12544 6507 12571 6534
rect 9305 6455 9331 6481
rect 9631 6453 9658 6480
rect 9916 6455 9942 6481
rect 10239 6453 10266 6480
rect 10527 6455 10553 6481
rect 10850 6453 10877 6480
rect 11105 6455 11131 6481
rect 11431 6453 11458 6480
rect 11716 6455 11742 6481
rect 12039 6453 12066 6480
rect 12327 6455 12353 6481
rect 12650 6453 12677 6480
rect 9405 6401 9431 6427
rect 9775 6417 9801 6443
rect 10016 6401 10042 6427
rect 10386 6417 10412 6443
rect 10627 6401 10653 6427
rect 10997 6417 11023 6443
rect 11205 6401 11231 6427
rect 11575 6417 11601 6443
rect 11816 6401 11842 6427
rect 12186 6417 12212 6443
rect 12427 6401 12453 6427
rect 12797 6417 12823 6443
rect 9521 5857 9548 5884
rect 11321 5857 11348 5884
rect 9305 5805 9331 5831
rect 9631 5803 9658 5830
rect 9916 5805 9942 5831
rect 10527 5805 10553 5831
rect 11105 5805 11131 5831
rect 11431 5803 11458 5830
rect 11716 5805 11742 5831
rect 12327 5805 12353 5831
rect 9405 5751 9431 5777
rect 9775 5767 9801 5793
rect 10016 5751 10042 5777
rect 10386 5767 10412 5793
rect 10627 5751 10653 5777
rect 10997 5767 11023 5793
rect 11205 5751 11231 5777
rect 11575 5767 11601 5793
rect 11816 5751 11842 5777
rect 12186 5767 12212 5793
rect 12427 5751 12453 5777
rect 12797 5767 12823 5793
rect 9519 5207 9546 5234
rect 10133 5206 10160 5233
rect 10743 5206 10770 5233
rect 11319 5207 11346 5234
rect 11933 5206 11960 5233
rect 12543 5206 12570 5233
rect 9305 5155 9331 5181
rect 9631 5153 9658 5180
rect 9916 5155 9942 5181
rect 10239 5153 10266 5180
rect 10527 5155 10553 5181
rect 10851 5153 10878 5180
rect 11105 5155 11131 5181
rect 11431 5153 11458 5180
rect 11716 5155 11742 5181
rect 12039 5153 12066 5180
rect 12327 5155 12353 5181
rect 12651 5153 12678 5180
rect 9405 5101 9431 5127
rect 9775 5117 9801 5143
rect 10016 5101 10042 5127
rect 10386 5117 10412 5143
rect 10627 5101 10653 5127
rect 10997 5117 11023 5143
rect 11205 5101 11231 5127
rect 11575 5117 11601 5143
rect 11816 5101 11842 5127
rect 12186 5117 12212 5143
rect 12427 5101 12453 5127
rect 12797 5117 12823 5143
rect 9519 4567 9546 4594
rect 10133 4567 10160 4594
rect 10744 4567 10771 4594
rect 11319 4567 11346 4594
rect 11933 4567 11960 4594
rect 12544 4567 12571 4594
rect 9305 4515 9331 4541
rect 9631 4513 9658 4540
rect 9916 4515 9942 4541
rect 10239 4513 10266 4540
rect 10527 4515 10553 4541
rect 10850 4513 10877 4540
rect 11105 4515 11131 4541
rect 11431 4513 11458 4540
rect 11716 4515 11742 4541
rect 12039 4513 12066 4540
rect 12327 4515 12353 4541
rect 12650 4513 12677 4540
rect 9405 4461 9431 4487
rect 9775 4477 9801 4503
rect 10016 4461 10042 4487
rect 10386 4477 10412 4503
rect 10627 4461 10653 4487
rect 10997 4477 11023 4503
rect 11205 4461 11231 4487
rect 11575 4477 11601 4503
rect 11816 4461 11842 4487
rect 12186 4477 12212 4503
rect 12427 4461 12453 4487
rect 12797 4477 12823 4503
rect 154 1113 186 1145
rect 13274 850 13314 890
rect 15206 850 15246 890
<< metal2 >>
rect 9302 7771 9335 8136
rect 9302 7745 9305 7771
rect 9331 7745 9335 7771
rect 9302 7121 9335 7745
rect 9302 7095 9305 7121
rect 9331 7095 9335 7121
rect 9302 6481 9335 7095
rect 9302 6455 9305 6481
rect 9331 6455 9335 6481
rect 9302 5831 9335 6455
rect 9302 5805 9305 5831
rect 9331 5805 9335 5831
rect 9302 5181 9335 5805
rect 9302 5155 9305 5181
rect 9331 5155 9335 5181
rect 9302 4541 9335 5155
rect 9302 4515 9305 4541
rect 9331 4515 9335 4541
rect 9302 4247 9335 4515
rect 9402 7717 9435 8136
rect 9402 7691 9405 7717
rect 9431 7691 9435 7717
rect 9402 7067 9435 7691
rect 9518 7824 9553 8136
rect 9518 7797 9521 7824
rect 9548 7797 9553 7824
rect 9518 7177 9553 7797
rect 9516 7174 9553 7177
rect 9516 7147 9519 7174
rect 9546 7147 9553 7174
rect 9516 7144 9553 7147
rect 9402 7041 9405 7067
rect 9431 7041 9435 7067
rect 9402 6427 9435 7041
rect 9518 6537 9553 7144
rect 9402 6401 9405 6427
rect 9431 6401 9435 6427
rect 9402 5777 9435 6401
rect 9516 6534 9553 6537
rect 9516 6507 9519 6534
rect 9546 6507 9553 6534
rect 9516 6188 9553 6507
rect 9402 5751 9405 5777
rect 9431 5751 9435 5777
rect 9402 5127 9435 5751
rect 9518 5884 9553 6188
rect 9518 5857 9521 5884
rect 9548 5857 9553 5884
rect 9518 5237 9553 5857
rect 9516 5234 9553 5237
rect 9516 5207 9519 5234
rect 9546 5207 9553 5234
rect 9516 5204 9553 5207
rect 9402 5101 9405 5127
rect 9431 5101 9435 5127
rect 9402 4487 9435 5101
rect 9518 4597 9553 5204
rect 9402 4461 9405 4487
rect 9431 4461 9435 4487
rect 9402 4247 9435 4461
rect 9516 4594 9553 4597
rect 9516 4567 9519 4594
rect 9546 4567 9553 4594
rect 9516 4248 9553 4567
rect 9624 7770 9661 8136
rect 9624 7743 9631 7770
rect 9658 7743 9661 7770
rect 9624 7120 9661 7743
rect 9624 7093 9631 7120
rect 9658 7093 9661 7120
rect 9624 6480 9661 7093
rect 9624 6453 9631 6480
rect 9658 6453 9661 6480
rect 9624 5830 9661 6453
rect 9624 5803 9631 5830
rect 9658 5803 9661 5830
rect 9624 5180 9661 5803
rect 9624 5153 9631 5180
rect 9658 5153 9661 5180
rect 9624 4540 9661 5153
rect 9624 4513 9631 4540
rect 9658 4513 9661 4540
rect 9624 4245 9661 4513
rect 9772 7733 9805 8136
rect 9772 7707 9775 7733
rect 9801 7707 9805 7733
rect 9772 7083 9805 7707
rect 9772 7057 9775 7083
rect 9801 7057 9805 7083
rect 9772 6443 9805 7057
rect 9772 6417 9775 6443
rect 9801 6417 9805 6443
rect 9772 5793 9805 6417
rect 9772 5767 9775 5793
rect 9801 5767 9805 5793
rect 9772 5143 9805 5767
rect 9772 5117 9775 5143
rect 9801 5117 9805 5143
rect 9772 4503 9805 5117
rect 9772 4477 9775 4503
rect 9801 4477 9805 4503
rect 9772 4247 9805 4477
rect 9913 7771 9946 8136
rect 9913 7745 9916 7771
rect 9942 7745 9946 7771
rect 9913 7121 9946 7745
rect 9913 7095 9916 7121
rect 9942 7095 9946 7121
rect 9913 6481 9946 7095
rect 9913 6455 9916 6481
rect 9942 6455 9946 6481
rect 9913 5831 9946 6455
rect 9913 5805 9916 5831
rect 9942 5805 9946 5831
rect 9913 5181 9946 5805
rect 9913 5155 9916 5181
rect 9942 5155 9946 5181
rect 9913 4541 9946 5155
rect 9913 4515 9916 4541
rect 9942 4515 9946 4541
rect 9913 4247 9946 4515
rect 10013 7717 10046 8136
rect 10013 7691 10016 7717
rect 10042 7691 10046 7717
rect 10013 7067 10046 7691
rect 10013 7041 10016 7067
rect 10042 7041 10046 7067
rect 10013 6427 10046 7041
rect 10013 6401 10016 6427
rect 10042 6401 10046 6427
rect 10013 5777 10046 6401
rect 10013 5751 10016 5777
rect 10042 5751 10046 5777
rect 10013 5127 10046 5751
rect 10013 5101 10016 5127
rect 10042 5101 10046 5127
rect 10013 4487 10046 5101
rect 10013 4461 10016 4487
rect 10042 4461 10046 4487
rect 10013 4247 10046 4461
rect 10127 7173 10164 8136
rect 10127 7146 10133 7173
rect 10160 7146 10164 7173
rect 10127 6534 10164 7146
rect 10127 6507 10133 6534
rect 10160 6507 10164 6534
rect 10127 5233 10164 6507
rect 10127 5206 10133 5233
rect 10160 5206 10164 5233
rect 10127 4594 10164 5206
rect 10127 4567 10133 4594
rect 10160 4567 10164 4594
rect 10127 4250 10164 4567
rect 10235 7120 10272 8136
rect 10235 7093 10239 7120
rect 10266 7093 10272 7120
rect 10235 6480 10272 7093
rect 10235 6453 10239 6480
rect 10266 6453 10272 6480
rect 10235 5180 10272 6453
rect 10235 5153 10239 5180
rect 10266 5153 10272 5180
rect 10235 4540 10272 5153
rect 10235 4513 10239 4540
rect 10266 4513 10272 4540
rect 10235 4253 10272 4513
rect 10383 7733 10416 8136
rect 10383 7707 10386 7733
rect 10412 7707 10416 7733
rect 10383 7083 10416 7707
rect 10383 7057 10386 7083
rect 10412 7057 10416 7083
rect 10383 6443 10416 7057
rect 10383 6417 10386 6443
rect 10412 6417 10416 6443
rect 10383 5793 10416 6417
rect 10383 5767 10386 5793
rect 10412 5767 10416 5793
rect 10383 5143 10416 5767
rect 10383 5117 10386 5143
rect 10412 5117 10416 5143
rect 10383 4503 10416 5117
rect 10383 4477 10386 4503
rect 10412 4477 10416 4503
rect 10383 4247 10416 4477
rect 10524 7771 10557 8136
rect 10524 7745 10527 7771
rect 10553 7745 10557 7771
rect 10524 7121 10557 7745
rect 10524 7095 10527 7121
rect 10553 7095 10557 7121
rect 10524 6481 10557 7095
rect 10524 6455 10527 6481
rect 10553 6455 10557 6481
rect 10524 5831 10557 6455
rect 10524 5805 10527 5831
rect 10553 5805 10557 5831
rect 10524 5181 10557 5805
rect 10524 5155 10527 5181
rect 10553 5155 10557 5181
rect 10524 4541 10557 5155
rect 10524 4515 10527 4541
rect 10553 4515 10557 4541
rect 10524 4247 10557 4515
rect 10624 7717 10657 8136
rect 10624 7691 10627 7717
rect 10653 7691 10657 7717
rect 10624 7067 10657 7691
rect 10624 7041 10627 7067
rect 10653 7041 10657 7067
rect 10624 6427 10657 7041
rect 10624 6401 10627 6427
rect 10653 6401 10657 6427
rect 10624 5777 10657 6401
rect 10624 5751 10627 5777
rect 10653 5751 10657 5777
rect 10624 5127 10657 5751
rect 10624 5101 10627 5127
rect 10653 5101 10657 5127
rect 10624 4487 10657 5101
rect 10624 4461 10627 4487
rect 10653 4461 10657 4487
rect 10624 4247 10657 4461
rect 10738 7173 10775 8136
rect 10738 7146 10743 7173
rect 10770 7146 10775 7173
rect 10738 6534 10775 7146
rect 10738 6507 10744 6534
rect 10771 6507 10775 6534
rect 10738 5233 10775 6507
rect 10738 5206 10743 5233
rect 10770 5206 10775 5233
rect 10738 4594 10775 5206
rect 10738 4567 10744 4594
rect 10771 4567 10775 4594
rect 10738 4251 10775 4567
rect 10846 7120 10883 8136
rect 10846 7093 10851 7120
rect 10878 7093 10883 7120
rect 10846 6480 10883 7093
rect 10846 6453 10850 6480
rect 10877 6453 10883 6480
rect 10846 5180 10883 6453
rect 10846 5153 10851 5180
rect 10878 5153 10883 5180
rect 10846 4540 10883 5153
rect 10846 4513 10850 4540
rect 10877 4513 10883 4540
rect 10846 4252 10883 4513
rect 10994 7733 11027 8136
rect 10994 7707 10997 7733
rect 11023 7707 11027 7733
rect 10994 7083 11027 7707
rect 10994 7057 10997 7083
rect 11023 7057 11027 7083
rect 10994 6443 11027 7057
rect 10994 6417 10997 6443
rect 11023 6417 11027 6443
rect 10994 5793 11027 6417
rect 10994 5767 10997 5793
rect 11023 5767 11027 5793
rect 10994 5143 11027 5767
rect 10994 5117 10997 5143
rect 11023 5117 11027 5143
rect 10994 4503 11027 5117
rect 10994 4477 10997 4503
rect 11023 4477 11027 4503
rect 10994 4247 11027 4477
rect 11102 7771 11135 8136
rect 11102 7745 11105 7771
rect 11131 7745 11135 7771
rect 11102 7121 11135 7745
rect 11102 7095 11105 7121
rect 11131 7095 11135 7121
rect 11102 6481 11135 7095
rect 11102 6455 11105 6481
rect 11131 6455 11135 6481
rect 11102 5831 11135 6455
rect 11102 5805 11105 5831
rect 11131 5805 11135 5831
rect 11102 5181 11135 5805
rect 11102 5155 11105 5181
rect 11131 5155 11135 5181
rect 11102 4541 11135 5155
rect 11102 4515 11105 4541
rect 11131 4515 11135 4541
rect 11102 4247 11135 4515
rect 11202 7717 11235 8136
rect 11202 7691 11205 7717
rect 11231 7691 11235 7717
rect 11202 7067 11235 7691
rect 11318 7824 11353 8136
rect 11318 7797 11321 7824
rect 11348 7797 11353 7824
rect 11318 7177 11353 7797
rect 11316 7174 11353 7177
rect 11316 7147 11319 7174
rect 11346 7147 11353 7174
rect 11316 7144 11353 7147
rect 11202 7041 11205 7067
rect 11231 7041 11235 7067
rect 11202 6427 11235 7041
rect 11318 6537 11353 7144
rect 11202 6401 11205 6427
rect 11231 6401 11235 6427
rect 11202 5777 11235 6401
rect 11316 6534 11353 6537
rect 11316 6507 11319 6534
rect 11346 6507 11353 6534
rect 11316 6188 11353 6507
rect 11202 5751 11205 5777
rect 11231 5751 11235 5777
rect 11202 5127 11235 5751
rect 11318 5884 11353 6188
rect 11318 5857 11321 5884
rect 11348 5857 11353 5884
rect 11318 5237 11353 5857
rect 11316 5234 11353 5237
rect 11316 5207 11319 5234
rect 11346 5207 11353 5234
rect 11316 5204 11353 5207
rect 11202 5101 11205 5127
rect 11231 5101 11235 5127
rect 11202 4487 11235 5101
rect 11318 4597 11353 5204
rect 11202 4461 11205 4487
rect 11231 4461 11235 4487
rect 11202 4247 11235 4461
rect 11316 4594 11353 4597
rect 11316 4567 11319 4594
rect 11346 4567 11353 4594
rect 11316 4248 11353 4567
rect 11424 7770 11461 8136
rect 11424 7743 11431 7770
rect 11458 7743 11461 7770
rect 11424 7120 11461 7743
rect 11424 7093 11431 7120
rect 11458 7093 11461 7120
rect 11424 6480 11461 7093
rect 11424 6453 11431 6480
rect 11458 6453 11461 6480
rect 11424 5830 11461 6453
rect 11424 5803 11431 5830
rect 11458 5803 11461 5830
rect 11424 5180 11461 5803
rect 11424 5153 11431 5180
rect 11458 5153 11461 5180
rect 11424 4540 11461 5153
rect 11424 4513 11431 4540
rect 11458 4513 11461 4540
rect 11424 4245 11461 4513
rect 11572 7733 11605 8136
rect 11572 7707 11575 7733
rect 11601 7707 11605 7733
rect 11572 7083 11605 7707
rect 11572 7057 11575 7083
rect 11601 7057 11605 7083
rect 11572 6443 11605 7057
rect 11572 6417 11575 6443
rect 11601 6417 11605 6443
rect 11572 5793 11605 6417
rect 11572 5767 11575 5793
rect 11601 5767 11605 5793
rect 11572 5143 11605 5767
rect 11572 5117 11575 5143
rect 11601 5117 11605 5143
rect 11572 4503 11605 5117
rect 11572 4477 11575 4503
rect 11601 4477 11605 4503
rect 11572 4247 11605 4477
rect 11713 7771 11746 8136
rect 11713 7745 11716 7771
rect 11742 7745 11746 7771
rect 11713 7121 11746 7745
rect 11713 7095 11716 7121
rect 11742 7095 11746 7121
rect 11713 6481 11746 7095
rect 11713 6455 11716 6481
rect 11742 6455 11746 6481
rect 11713 5831 11746 6455
rect 11713 5805 11716 5831
rect 11742 5805 11746 5831
rect 11713 5181 11746 5805
rect 11713 5155 11716 5181
rect 11742 5155 11746 5181
rect 11713 4541 11746 5155
rect 11713 4515 11716 4541
rect 11742 4515 11746 4541
rect 11713 4247 11746 4515
rect 11813 7717 11846 8136
rect 11813 7691 11816 7717
rect 11842 7691 11846 7717
rect 11813 7067 11846 7691
rect 11813 7041 11816 7067
rect 11842 7041 11846 7067
rect 11813 6427 11846 7041
rect 11813 6401 11816 6427
rect 11842 6401 11846 6427
rect 11813 5777 11846 6401
rect 11813 5751 11816 5777
rect 11842 5751 11846 5777
rect 11813 5127 11846 5751
rect 11813 5101 11816 5127
rect 11842 5101 11846 5127
rect 11813 4487 11846 5101
rect 11813 4461 11816 4487
rect 11842 4461 11846 4487
rect 11813 4247 11846 4461
rect 11927 7173 11964 8136
rect 11927 7146 11933 7173
rect 11960 7146 11964 7173
rect 11927 6534 11964 7146
rect 11927 6507 11933 6534
rect 11960 6507 11964 6534
rect 11927 5233 11964 6507
rect 11927 5206 11933 5233
rect 11960 5206 11964 5233
rect 11927 4594 11964 5206
rect 11927 4567 11933 4594
rect 11960 4567 11964 4594
rect 11927 4250 11964 4567
rect 12035 7120 12072 8136
rect 12035 7093 12039 7120
rect 12066 7093 12072 7120
rect 12035 6480 12072 7093
rect 12035 6453 12039 6480
rect 12066 6453 12072 6480
rect 12035 5180 12072 6453
rect 12035 5153 12039 5180
rect 12066 5153 12072 5180
rect 12035 4540 12072 5153
rect 12035 4513 12039 4540
rect 12066 4513 12072 4540
rect 12035 4253 12072 4513
rect 12183 7733 12216 8136
rect 12183 7707 12186 7733
rect 12212 7707 12216 7733
rect 12183 7083 12216 7707
rect 12183 7057 12186 7083
rect 12212 7057 12216 7083
rect 12183 6443 12216 7057
rect 12183 6417 12186 6443
rect 12212 6417 12216 6443
rect 12183 5793 12216 6417
rect 12183 5767 12186 5793
rect 12212 5767 12216 5793
rect 12183 5143 12216 5767
rect 12183 5117 12186 5143
rect 12212 5117 12216 5143
rect 12183 4503 12216 5117
rect 12183 4477 12186 4503
rect 12212 4477 12216 4503
rect 12183 4247 12216 4477
rect 12324 7771 12357 8136
rect 12324 7745 12327 7771
rect 12353 7745 12357 7771
rect 12324 7121 12357 7745
rect 12324 7095 12327 7121
rect 12353 7095 12357 7121
rect 12324 6481 12357 7095
rect 12324 6455 12327 6481
rect 12353 6455 12357 6481
rect 12324 5831 12357 6455
rect 12324 5805 12327 5831
rect 12353 5805 12357 5831
rect 12324 5181 12357 5805
rect 12324 5155 12327 5181
rect 12353 5155 12357 5181
rect 12324 4541 12357 5155
rect 12324 4515 12327 4541
rect 12353 4515 12357 4541
rect 12324 4247 12357 4515
rect 12424 7717 12457 8136
rect 12424 7691 12427 7717
rect 12453 7691 12457 7717
rect 12424 7067 12457 7691
rect 12424 7041 12427 7067
rect 12453 7041 12457 7067
rect 12424 6427 12457 7041
rect 12424 6401 12427 6427
rect 12453 6401 12457 6427
rect 12424 5777 12457 6401
rect 12424 5751 12427 5777
rect 12453 5751 12457 5777
rect 12424 5127 12457 5751
rect 12424 5101 12427 5127
rect 12453 5101 12457 5127
rect 12424 4487 12457 5101
rect 12424 4461 12427 4487
rect 12453 4461 12457 4487
rect 12424 4247 12457 4461
rect 12538 7173 12575 8136
rect 12538 7146 12543 7173
rect 12570 7146 12575 7173
rect 12538 6534 12575 7146
rect 12538 6507 12544 6534
rect 12571 6507 12575 6534
rect 12538 5233 12575 6507
rect 12538 5206 12543 5233
rect 12570 5206 12575 5233
rect 12538 4594 12575 5206
rect 12538 4567 12544 4594
rect 12571 4567 12575 4594
rect 12538 4251 12575 4567
rect 12646 7120 12683 8136
rect 12646 7093 12651 7120
rect 12678 7093 12683 7120
rect 12646 6480 12683 7093
rect 12646 6453 12650 6480
rect 12677 6453 12683 6480
rect 12646 5180 12683 6453
rect 12646 5153 12651 5180
rect 12678 5153 12683 5180
rect 12646 4540 12683 5153
rect 12646 4513 12650 4540
rect 12677 4513 12683 4540
rect 12646 4252 12683 4513
rect 12794 7733 12827 8136
rect 12794 7707 12797 7733
rect 12823 7707 12827 7733
rect 12794 7083 12827 7707
rect 12794 7057 12797 7083
rect 12823 7057 12827 7083
rect 12794 6443 12827 7057
rect 12794 6417 12797 6443
rect 12823 6417 12827 6443
rect 12794 5793 12827 6417
rect 12794 5767 12797 5793
rect 12823 5767 12827 5793
rect 12794 5143 12827 5767
rect 12794 5117 12797 5143
rect 12823 5117 12827 5143
rect 12794 4503 12827 5117
rect 12794 4477 12797 4503
rect 12823 4477 12827 4503
rect 12794 4247 12827 4477
rect 100 1145 300 1154
rect 100 1113 154 1145
rect 186 1113 300 1145
rect 100 1104 300 1113
rect 13249 890 13339 915
rect 13249 850 13274 890
rect 13314 850 13339 890
rect 13249 825 13339 850
rect 15181 890 15271 915
rect 15181 850 15206 890
rect 15246 850 15271 890
rect 15181 825 15271 850
rect 400 674 600 683
rect 400 642 466 674
rect 498 642 600 674
rect 400 633 600 642
<< via2 >>
rect 154 1113 186 1145
rect 13274 850 13314 890
rect 15206 850 15246 890
rect 466 642 498 674
<< metal3 >>
rect 100 1145 300 1154
rect 100 1113 154 1145
rect 186 1113 300 1145
rect 100 1104 300 1113
rect 13249 890 13339 915
rect 13249 850 13274 890
rect 13314 850 13339 890
rect 13249 825 13339 850
rect 15181 890 15271 915
rect 15181 850 15206 890
rect 15246 850 15271 890
rect 15181 825 15271 850
rect 400 674 600 683
rect 400 642 466 674
rect 498 642 600 674
rect 400 633 600 642
<< via3 >>
rect 154 1113 186 1145
rect 13274 850 13314 890
rect 15206 850 15246 890
rect 466 642 498 674
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 7483 22476 7513 22576
rect 7759 22476 7789 22576
rect 8035 22476 8065 22576
rect 8311 22476 8341 22576
rect 8587 22476 8617 22576
rect 8863 22476 8893 22576
rect 9139 22476 9169 22576
rect 9415 22476 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 100 1145 300 22076
rect 100 1113 154 1145
rect 186 1113 300 1145
rect 100 500 300 1113
rect 400 674 600 22076
rect 400 642 466 674
rect 498 642 600 674
rect 400 500 600 642
rect 13249 890 13339 915
rect 13249 850 13274 890
rect 13314 850 13339 890
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 850
rect 15181 890 15271 915
rect 15181 850 15206 890
rect 15246 850 15271 890
rect 15181 0 15271 850
use latch_sr  latch_sr_0
timestamp 1753205587
transform 1 0 9452 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_1
timestamp 1753205587
transform 1 0 9452 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_2
timestamp 1753205587
transform 1 0 9452 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_3
timestamp 1753205587
transform 1 0 10063 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_4
timestamp 1753205587
transform 1 0 10063 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_5
timestamp 1753205587
transform 1 0 10063 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_6
timestamp 1753205587
transform 1 0 10674 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_7
timestamp 1753205587
transform 1 0 10674 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_8
timestamp 1753205587
transform 1 0 10674 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_9
timestamp 1753205587
transform 1 0 11252 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_10
timestamp 1753205587
transform 1 0 11863 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_11
timestamp 1753205587
transform 1 0 12474 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_12
timestamp 1753205587
transform 1 0 11252 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_13
timestamp 1753205587
transform 1 0 11863 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_14
timestamp 1753205587
transform 1 0 12474 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_15
timestamp 1753205587
transform 1 0 11252 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_16
timestamp 1753205587
transform 1 0 11863 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_17
timestamp 1753205587
transform 1 0 12474 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_18
timestamp 1753205587
transform 1 0 12474 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_19
timestamp 1753205587
transform 1 0 11863 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_20
timestamp 1753205587
transform 1 0 11252 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_21
timestamp 1753205587
transform 1 0 10674 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_22
timestamp 1753205587
transform 1 0 10063 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_23
timestamp 1753205587
transform 1 0 9452 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_24
timestamp 1753205587
transform 1 0 12474 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_25
timestamp 1753205587
transform 1 0 11863 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_26
timestamp 1753205587
transform 1 0 11252 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_27
timestamp 1753205587
transform 1 0 10674 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_28
timestamp 1753205587
transform 1 0 10063 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_29
timestamp 1753205587
transform 1 0 9452 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_30
timestamp 1753205587
transform 1 0 12474 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_31
timestamp 1753205587
transform 1 0 11863 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_32
timestamp 1753205587
transform 1 0 11252 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_33
timestamp 1753205587
transform 1 0 10674 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_34
timestamp 1753205587
transform 1 0 10063 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_35
timestamp 1753205587
transform 1 0 9452 0 1 4340
box -2 -49 275 526
use NOT  NOT_0
timestamp 1750779130
transform 1 0 14171 0 1 657
box -87 -24 160 609
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
