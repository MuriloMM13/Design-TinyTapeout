VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOT
  CLASS CORE ;
  FOREIGN NOT ;
  ORIGIN 0.190 0.240 ;
  SIZE 1.790 BY 3.200 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT -0.190 1.080 0.630 1.280 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.442800 ;
    PORT
      LAYER li1 ;
        RECT 0.720 1.490 1.060 2.460 ;
        RECT 0.810 1.280 1.060 1.490 ;
        RECT 0.810 1.080 1.600 1.280 ;
        RECT 0.810 0.890 1.060 1.080 ;
        RECT 0.720 0.260 1.060 0.890 ;
    END
  END Y
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.310 1.490 0.540 2.630 ;
      LAYER met1 ;
        RECT -0.190 2.480 1.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.310 0.090 0.540 0.910 ;
        RECT 0.000 -0.090 1.380 0.090 ;
      LAYER met1 ;
        RECT -0.190 -0.240 1.600 0.240 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT -0.190 1.300 1.600 2.910 ;
      LAYER pwell ;
        RECT 0.210 0.910 0.720 1.020 ;
        RECT 0.210 0.890 0.550 0.910 ;
        RECT 0.560 0.890 0.720 0.910 ;
        RECT 0.810 0.890 1.140 1.020 ;
        RECT 0.210 -0.090 1.140 0.890 ;
  END
END NOT
END LIBRARY

