VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOT
  CLASS CORE ;
  FOREIGN NOT ;
  ORIGIN 0.810 0.240 ;
  SIZE 2.410 BY 3.200 ;
  SITE unithd ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT -0.290 2.480 0.140 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.290 -0.240 0.140 0.240 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT -0.810 1.090 -0.630 1.270 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.442800 ;
    PORT
      LAYER li1 ;
        RECT 0.810 1.080 1.600 1.280 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT -0.460 -0.160 1.600 2.910 ;
      LAYER li1 ;
        RECT -0.810 1.450 1.380 2.810 ;
        RECT -0.810 1.440 0.640 1.450 ;
        RECT -0.460 1.280 0.640 1.440 ;
        RECT -0.810 1.270 0.640 1.280 ;
        RECT -0.460 1.090 0.640 1.270 ;
        RECT -0.810 1.080 0.640 1.090 ;
        RECT -0.460 0.920 0.640 1.080 ;
        RECT -0.810 0.910 0.640 0.920 ;
        RECT -0.810 -0.090 1.380 0.910 ;
      LAYER met1 ;
        RECT 0.420 2.200 1.600 2.960 ;
        RECT 0.140 0.520 1.600 2.200 ;
        RECT 0.420 -0.240 1.600 0.520 ;
  END
END NOT
END LIBRARY

