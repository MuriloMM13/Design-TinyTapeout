VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOT
  CLASS CORE ;
  FOREIGN NOT ;
  ORIGIN 1.070 0.440 ;
  SIZE 2.870 BY 3.600 ;
  SITE unithd ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT -0.870 2.630 -0.690 2.810 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT -0.870 -0.090 -0.690 0.090 ;
    END
  END VGND
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT -0.870 1.090 -0.690 1.270 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.442800 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.090 1.600 1.270 ;
    END
  END Y
  OBS
      LAYER nwell ;
        RECT -0.870 1.290 1.600 2.910 ;
      LAYER pwell ;
        RECT -0.870 -0.190 1.600 1.020 ;
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.310 1.870 0.540 2.630 ;
        RECT -0.160 1.490 0.540 1.870 ;
        RECT 0.720 1.490 1.060 2.460 ;
        RECT 0.810 1.280 1.060 1.490 ;
        RECT -0.870 1.270 -0.500 1.280 ;
        RECT -0.690 1.090 -0.500 1.270 ;
        RECT -0.870 1.080 -0.500 1.090 ;
        RECT 0.810 1.270 1.600 1.280 ;
        RECT 0.810 1.090 1.420 1.270 ;
        RECT 0.810 1.080 1.600 1.090 ;
        RECT -0.330 0.550 0.540 0.910 ;
        RECT 0.810 0.890 1.060 1.080 ;
        RECT 0.310 0.090 0.540 0.550 ;
        RECT 0.720 0.260 1.060 0.890 ;
        RECT 0.000 -0.090 1.380 0.090 ;
      LAYER met1 ;
        RECT -0.870 2.810 1.600 2.960 ;
        RECT -0.690 2.630 1.600 2.810 ;
        RECT -0.870 2.480 1.600 2.630 ;
        RECT -0.870 0.090 1.600 0.240 ;
        RECT -0.690 -0.090 1.600 0.090 ;
        RECT -0.870 -0.240 1.600 -0.090 ;
  END
END NOT
END LIBRARY

