magic
tech sky130A
timestamp 1753205587
<< nwell >>
rect 50 256 223 492
<< nmos >>
rect 27 0 42 100
rect 63 0 78 100
rect 107 0 122 100
rect 151 0 166 100
rect 195 0 210 100
rect 231 0 246 100
<< pmos >>
rect 107 274 122 474
rect 151 274 166 474
<< ndiff >>
rect -2 93 27 100
rect -2 76 4 93
rect 21 76 27 93
rect -2 59 27 76
rect -2 42 4 59
rect 21 42 27 59
rect -2 25 27 42
rect -2 8 4 25
rect 21 8 27 25
rect -2 0 27 8
rect 42 0 63 100
rect 78 93 107 100
rect 78 76 84 93
rect 101 76 107 93
rect 78 59 107 76
rect 78 42 84 59
rect 101 42 107 59
rect 78 25 107 42
rect 78 8 84 25
rect 101 8 107 25
rect 78 0 107 8
rect 122 93 151 100
rect 122 76 128 93
rect 145 76 151 93
rect 122 59 151 76
rect 122 42 128 59
rect 145 42 151 59
rect 122 25 151 42
rect 122 8 128 25
rect 145 8 151 25
rect 122 0 151 8
rect 166 93 195 100
rect 166 76 172 93
rect 189 76 195 93
rect 166 59 195 76
rect 166 42 172 59
rect 189 42 195 59
rect 166 25 195 42
rect 166 8 172 25
rect 189 8 195 25
rect 166 0 195 8
rect 210 0 231 100
rect 246 93 275 100
rect 246 76 252 93
rect 269 76 275 93
rect 246 59 275 76
rect 246 42 252 59
rect 269 42 275 59
rect 246 25 275 42
rect 246 8 252 25
rect 269 8 275 25
rect 246 0 275 8
<< pdiff >>
rect 78 469 107 474
rect 78 452 84 469
rect 101 452 107 469
rect 78 435 107 452
rect 78 418 84 435
rect 101 418 107 435
rect 78 401 107 418
rect 78 384 84 401
rect 101 384 107 401
rect 78 367 107 384
rect 78 350 84 367
rect 101 350 107 367
rect 78 333 107 350
rect 78 316 84 333
rect 101 316 107 333
rect 78 299 107 316
rect 78 282 84 299
rect 101 282 107 299
rect 78 274 107 282
rect 122 469 151 474
rect 122 452 128 469
rect 145 452 151 469
rect 122 435 151 452
rect 122 418 128 435
rect 145 418 151 435
rect 122 401 151 418
rect 122 384 128 401
rect 145 384 151 401
rect 122 367 151 384
rect 122 350 128 367
rect 145 350 151 367
rect 122 333 151 350
rect 122 316 128 333
rect 145 316 151 333
rect 122 299 151 316
rect 122 282 128 299
rect 145 282 151 299
rect 122 274 151 282
rect 166 469 195 474
rect 166 452 172 469
rect 189 452 195 469
rect 166 435 195 452
rect 166 418 172 435
rect 189 418 195 435
rect 166 401 195 418
rect 166 384 172 401
rect 189 384 195 401
rect 166 367 195 384
rect 166 350 172 367
rect 189 350 195 367
rect 166 333 195 350
rect 166 316 172 333
rect 189 316 195 333
rect 166 299 195 316
rect 166 282 172 299
rect 189 282 195 299
rect 166 274 195 282
<< ndiffc >>
rect 4 76 21 93
rect 4 42 21 59
rect 4 8 21 25
rect 84 76 101 93
rect 84 42 101 59
rect 84 8 101 25
rect 128 76 145 93
rect 128 42 145 59
rect 128 8 145 25
rect 172 76 189 93
rect 172 42 189 59
rect 172 8 189 25
rect 252 76 269 93
rect 252 42 269 59
rect 252 8 269 25
<< pdiffc >>
rect 84 452 101 469
rect 84 418 101 435
rect 84 384 101 401
rect 84 350 101 367
rect 84 316 101 333
rect 84 282 101 299
rect 128 452 145 469
rect 128 418 145 435
rect 128 384 145 401
rect 128 350 145 367
rect 128 316 145 333
rect 128 282 145 299
rect 172 452 189 469
rect 172 418 189 435
rect 172 384 189 401
rect 172 350 189 367
rect 172 316 189 333
rect 172 282 189 299
<< poly >>
rect 107 474 122 487
rect 151 474 166 487
rect 107 257 122 274
rect 97 249 130 257
rect 97 232 105 249
rect 122 232 130 249
rect 97 224 130 232
rect -2 197 31 205
rect -2 180 6 197
rect 23 187 31 197
rect 23 180 78 187
rect -2 172 78 180
rect -2 143 42 151
rect -2 126 6 143
rect 23 126 42 143
rect -2 118 42 126
rect 27 100 42 118
rect 63 100 78 172
rect 107 100 122 224
rect 151 203 166 274
rect 143 195 176 203
rect 143 178 151 195
rect 168 178 176 195
rect 143 170 176 178
rect 151 100 166 170
rect 242 159 275 167
rect 242 149 250 159
rect 195 142 250 149
rect 267 142 275 159
rect 195 134 275 142
rect 195 100 210 134
rect 231 100 246 113
rect 27 -34 42 0
rect 63 -13 78 0
rect 107 -13 122 0
rect 151 -13 166 0
rect 195 -13 210 0
rect 231 -34 246 0
rect 27 -49 246 -34
<< polycont >>
rect 105 232 122 249
rect 6 180 23 197
rect 6 126 23 143
rect 151 178 168 195
rect 250 142 267 159
<< locali >>
rect 123 492 127 511
rect 146 492 150 511
rect 48 469 106 477
rect 48 452 84 469
rect 101 452 106 469
rect 48 435 106 452
rect 48 418 84 435
rect 101 418 106 435
rect 48 401 106 418
rect 48 384 84 401
rect 101 384 106 401
rect 48 367 106 384
rect 48 350 84 367
rect 101 350 106 367
rect 48 333 106 350
rect 48 316 84 333
rect 101 316 106 333
rect 48 299 106 316
rect 48 282 84 299
rect 101 282 106 299
rect 48 274 106 282
rect 123 469 150 492
rect 123 452 128 469
rect 145 452 150 469
rect 123 435 150 452
rect 123 418 128 435
rect 145 418 150 435
rect 123 401 150 418
rect 123 384 128 401
rect 145 384 150 401
rect 123 367 150 384
rect 123 350 128 367
rect 145 350 150 367
rect 123 333 150 350
rect 123 316 128 333
rect 145 316 150 333
rect 123 299 150 316
rect 123 282 128 299
rect 145 282 150 299
rect 123 274 150 282
rect 167 469 225 477
rect 167 452 172 469
rect 189 452 225 469
rect 167 435 225 452
rect 167 418 172 435
rect 189 418 225 435
rect 167 401 225 418
rect 167 384 172 401
rect 189 384 225 401
rect 167 367 225 384
rect 167 350 172 367
rect 189 350 225 367
rect 167 333 225 350
rect 167 316 172 333
rect 189 316 225 333
rect 167 299 225 316
rect 167 282 172 299
rect 189 282 225 299
rect 167 274 225 282
rect -2 197 31 205
rect -2 180 6 197
rect 23 180 31 197
rect -2 172 31 180
rect 48 187 75 274
rect 97 249 130 257
rect 97 232 105 249
rect 122 241 130 249
rect 198 241 225 274
rect 122 232 225 241
rect 97 224 225 232
rect 143 195 176 203
rect 143 187 151 195
rect 48 178 151 187
rect 168 178 176 195
rect 48 170 176 178
rect -2 143 31 151
rect -2 126 6 143
rect 23 126 31 143
rect -2 118 31 126
rect 48 101 75 170
rect 198 101 225 224
rect 242 159 275 167
rect 242 142 250 159
rect 267 142 275 159
rect 242 134 275 142
rect -1 93 26 101
rect -1 76 4 93
rect 21 76 26 93
rect -1 59 26 76
rect -1 42 4 59
rect 21 42 26 59
rect -1 25 26 42
rect -1 8 4 25
rect 21 8 26 25
rect -1 0 26 8
rect 48 93 106 101
rect 48 76 84 93
rect 101 76 106 93
rect 48 59 106 76
rect 48 42 84 59
rect 101 42 106 59
rect 48 25 106 42
rect 48 8 84 25
rect 101 8 106 25
rect 48 0 106 8
rect 123 93 150 101
rect 123 76 128 93
rect 145 76 150 93
rect 123 59 150 76
rect 123 42 128 59
rect 145 42 150 59
rect 123 25 150 42
rect 123 8 128 25
rect 145 8 150 25
rect 123 -15 150 8
rect 167 93 225 101
rect 167 76 172 93
rect 189 76 225 93
rect 167 59 225 76
rect 167 42 172 59
rect 189 42 225 59
rect 167 25 225 42
rect 167 8 172 25
rect 189 8 225 25
rect 167 0 225 8
rect 247 93 274 101
rect 247 76 252 93
rect 269 76 274 93
rect 247 59 274 76
rect 247 42 252 59
rect 269 42 274 59
rect 247 25 274 42
rect 247 8 252 25
rect 269 8 274 25
rect 247 0 274 8
rect 123 -34 127 -15
rect 146 -34 150 -15
<< viali >>
rect 127 492 146 511
rect 6 180 23 197
rect 105 232 122 249
rect 151 178 168 195
rect 6 126 23 143
rect 250 142 267 159
rect 127 -34 146 -15
<< metal1 >>
rect -2 511 275 526
rect -2 492 127 511
rect 146 492 275 511
rect -2 477 275 492
rect 97 249 130 257
rect 97 232 105 249
rect 122 232 130 249
rect 97 224 130 232
rect -2 197 31 205
rect -2 180 6 197
rect 23 180 31 197
rect -2 172 31 180
rect 143 195 176 203
rect 143 178 151 195
rect 168 178 176 195
rect 143 170 176 178
rect 242 159 275 167
rect -2 143 31 151
rect -2 126 6 143
rect 23 126 31 143
rect 242 142 250 159
rect 267 142 275 159
rect 242 134 275 142
rect -2 118 31 126
rect -2 -15 275 0
rect -2 -34 127 -15
rect 146 -34 275 -15
rect -2 -49 275 -34
<< end >>
