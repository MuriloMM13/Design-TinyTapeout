* NGSPICE file created from tt_um_analog_murilo.ext - technology: sky130A

.subckt NOT VGND VDPWR A Y
X0 Y A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2673 pd=2.52 as=0.2673 ps=2.52 w=0.99 l=0.15
X1 Y A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.1755 ps=1.84 w=0.65 l=0.15
.ends

.subckt tt_um_analog_murilo clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
XNOT_0 SUB VDPWR ua[1] ua[0] NOT
.ends

