magic
tech sky130A
timestamp 1753208296
<< nwell >>
rect 13113 7826 13286 8062
rect 13724 7826 13897 8062
rect 14302 7826 14475 8062
rect 14913 7826 15086 8062
rect 15524 7826 15697 8062
rect 12502 7176 12675 7412
rect 13113 7176 13286 7412
rect 13724 7176 13897 7412
rect 14302 7176 14475 7412
rect 14913 7176 15086 7412
rect 15524 7176 15697 7412
rect 12502 6536 12675 6772
rect 13113 6536 13286 6772
rect 13724 6536 13897 6772
rect 14302 6536 14475 6772
rect 14913 6536 15086 6772
rect 15524 6536 15697 6772
rect 12502 5886 12675 6122
rect 13113 5886 13286 6122
rect 13724 5886 13897 6122
rect 14302 5886 14475 6122
rect 14913 5886 15086 6122
rect 15524 5886 15697 6122
rect 12502 5236 12675 5472
rect 13113 5236 13286 5472
rect 13724 5236 13897 5472
rect 14302 5236 14475 5472
rect 14913 5236 15086 5472
rect 15524 5236 15697 5472
rect 12502 4596 12675 4832
rect 13113 4596 13286 4832
rect 13724 4596 13897 4832
rect 14302 4596 14475 4832
rect 14913 4596 15086 4832
rect 15524 4596 15697 4832
<< nmos >>
rect 13090 7570 13105 7670
rect 13126 7570 13141 7670
rect 13170 7570 13185 7670
rect 13214 7570 13229 7670
rect 13258 7570 13273 7670
rect 13294 7570 13309 7670
rect 13701 7570 13716 7670
rect 13737 7570 13752 7670
rect 13781 7570 13796 7670
rect 13825 7570 13840 7670
rect 13869 7570 13884 7670
rect 13905 7570 13920 7670
rect 14279 7570 14294 7670
rect 14315 7570 14330 7670
rect 14359 7570 14374 7670
rect 14403 7570 14418 7670
rect 14447 7570 14462 7670
rect 14483 7570 14498 7670
rect 14890 7570 14905 7670
rect 14926 7570 14941 7670
rect 14970 7570 14985 7670
rect 15014 7570 15029 7670
rect 15058 7570 15073 7670
rect 15094 7570 15109 7670
rect 15501 7570 15516 7670
rect 15537 7570 15552 7670
rect 15581 7570 15596 7670
rect 15625 7570 15640 7670
rect 15669 7570 15684 7670
rect 15705 7570 15720 7670
rect 12479 6920 12494 7020
rect 12515 6920 12530 7020
rect 12559 6920 12574 7020
rect 12603 6920 12618 7020
rect 12647 6920 12662 7020
rect 12683 6920 12698 7020
rect 13090 6920 13105 7020
rect 13126 6920 13141 7020
rect 13170 6920 13185 7020
rect 13214 6920 13229 7020
rect 13258 6920 13273 7020
rect 13294 6920 13309 7020
rect 13701 6920 13716 7020
rect 13737 6920 13752 7020
rect 13781 6920 13796 7020
rect 13825 6920 13840 7020
rect 13869 6920 13884 7020
rect 13905 6920 13920 7020
rect 14279 6920 14294 7020
rect 14315 6920 14330 7020
rect 14359 6920 14374 7020
rect 14403 6920 14418 7020
rect 14447 6920 14462 7020
rect 14483 6920 14498 7020
rect 14890 6920 14905 7020
rect 14926 6920 14941 7020
rect 14970 6920 14985 7020
rect 15014 6920 15029 7020
rect 15058 6920 15073 7020
rect 15094 6920 15109 7020
rect 15501 6920 15516 7020
rect 15537 6920 15552 7020
rect 15581 6920 15596 7020
rect 15625 6920 15640 7020
rect 15669 6920 15684 7020
rect 15705 6920 15720 7020
rect 12479 6280 12494 6380
rect 12515 6280 12530 6380
rect 12559 6280 12574 6380
rect 12603 6280 12618 6380
rect 12647 6280 12662 6380
rect 12683 6280 12698 6380
rect 13090 6280 13105 6380
rect 13126 6280 13141 6380
rect 13170 6280 13185 6380
rect 13214 6280 13229 6380
rect 13258 6280 13273 6380
rect 13294 6280 13309 6380
rect 13701 6280 13716 6380
rect 13737 6280 13752 6380
rect 13781 6280 13796 6380
rect 13825 6280 13840 6380
rect 13869 6280 13884 6380
rect 13905 6280 13920 6380
rect 14279 6280 14294 6380
rect 14315 6280 14330 6380
rect 14359 6280 14374 6380
rect 14403 6280 14418 6380
rect 14447 6280 14462 6380
rect 14483 6280 14498 6380
rect 14890 6280 14905 6380
rect 14926 6280 14941 6380
rect 14970 6280 14985 6380
rect 15014 6280 15029 6380
rect 15058 6280 15073 6380
rect 15094 6280 15109 6380
rect 15501 6280 15516 6380
rect 15537 6280 15552 6380
rect 15581 6280 15596 6380
rect 15625 6280 15640 6380
rect 15669 6280 15684 6380
rect 15705 6280 15720 6380
rect 12479 5630 12494 5730
rect 12515 5630 12530 5730
rect 12559 5630 12574 5730
rect 12603 5630 12618 5730
rect 12647 5630 12662 5730
rect 12683 5630 12698 5730
rect 13090 5630 13105 5730
rect 13126 5630 13141 5730
rect 13170 5630 13185 5730
rect 13214 5630 13229 5730
rect 13258 5630 13273 5730
rect 13294 5630 13309 5730
rect 13701 5630 13716 5730
rect 13737 5630 13752 5730
rect 13781 5630 13796 5730
rect 13825 5630 13840 5730
rect 13869 5630 13884 5730
rect 13905 5630 13920 5730
rect 14279 5630 14294 5730
rect 14315 5630 14330 5730
rect 14359 5630 14374 5730
rect 14403 5630 14418 5730
rect 14447 5630 14462 5730
rect 14483 5630 14498 5730
rect 14890 5630 14905 5730
rect 14926 5630 14941 5730
rect 14970 5630 14985 5730
rect 15014 5630 15029 5730
rect 15058 5630 15073 5730
rect 15094 5630 15109 5730
rect 15501 5630 15516 5730
rect 15537 5630 15552 5730
rect 15581 5630 15596 5730
rect 15625 5630 15640 5730
rect 15669 5630 15684 5730
rect 15705 5630 15720 5730
rect 12479 4980 12494 5080
rect 12515 4980 12530 5080
rect 12559 4980 12574 5080
rect 12603 4980 12618 5080
rect 12647 4980 12662 5080
rect 12683 4980 12698 5080
rect 13090 4980 13105 5080
rect 13126 4980 13141 5080
rect 13170 4980 13185 5080
rect 13214 4980 13229 5080
rect 13258 4980 13273 5080
rect 13294 4980 13309 5080
rect 13701 4980 13716 5080
rect 13737 4980 13752 5080
rect 13781 4980 13796 5080
rect 13825 4980 13840 5080
rect 13869 4980 13884 5080
rect 13905 4980 13920 5080
rect 14279 4980 14294 5080
rect 14315 4980 14330 5080
rect 14359 4980 14374 5080
rect 14403 4980 14418 5080
rect 14447 4980 14462 5080
rect 14483 4980 14498 5080
rect 14890 4980 14905 5080
rect 14926 4980 14941 5080
rect 14970 4980 14985 5080
rect 15014 4980 15029 5080
rect 15058 4980 15073 5080
rect 15094 4980 15109 5080
rect 15501 4980 15516 5080
rect 15537 4980 15552 5080
rect 15581 4980 15596 5080
rect 15625 4980 15640 5080
rect 15669 4980 15684 5080
rect 15705 4980 15720 5080
rect 12479 4340 12494 4440
rect 12515 4340 12530 4440
rect 12559 4340 12574 4440
rect 12603 4340 12618 4440
rect 12647 4340 12662 4440
rect 12683 4340 12698 4440
rect 13090 4340 13105 4440
rect 13126 4340 13141 4440
rect 13170 4340 13185 4440
rect 13214 4340 13229 4440
rect 13258 4340 13273 4440
rect 13294 4340 13309 4440
rect 13701 4340 13716 4440
rect 13737 4340 13752 4440
rect 13781 4340 13796 4440
rect 13825 4340 13840 4440
rect 13869 4340 13884 4440
rect 13905 4340 13920 4440
rect 14279 4340 14294 4440
rect 14315 4340 14330 4440
rect 14359 4340 14374 4440
rect 14403 4340 14418 4440
rect 14447 4340 14462 4440
rect 14483 4340 14498 4440
rect 14890 4340 14905 4440
rect 14926 4340 14941 4440
rect 14970 4340 14985 4440
rect 15014 4340 15029 4440
rect 15058 4340 15073 4440
rect 15094 4340 15109 4440
rect 15501 4340 15516 4440
rect 15537 4340 15552 4440
rect 15581 4340 15596 4440
rect 15625 4340 15640 4440
rect 15669 4340 15684 4440
rect 15705 4340 15720 4440
<< pmos >>
rect 13170 7844 13185 8044
rect 13214 7844 13229 8044
rect 13781 7844 13796 8044
rect 13825 7844 13840 8044
rect 14359 7844 14374 8044
rect 14403 7844 14418 8044
rect 14970 7844 14985 8044
rect 15014 7844 15029 8044
rect 15581 7844 15596 8044
rect 15625 7844 15640 8044
rect 12559 7194 12574 7394
rect 12603 7194 12618 7394
rect 13170 7194 13185 7394
rect 13214 7194 13229 7394
rect 13781 7194 13796 7394
rect 13825 7194 13840 7394
rect 14359 7194 14374 7394
rect 14403 7194 14418 7394
rect 14970 7194 14985 7394
rect 15014 7194 15029 7394
rect 15581 7194 15596 7394
rect 15625 7194 15640 7394
rect 12559 6554 12574 6754
rect 12603 6554 12618 6754
rect 13170 6554 13185 6754
rect 13214 6554 13229 6754
rect 13781 6554 13796 6754
rect 13825 6554 13840 6754
rect 14359 6554 14374 6754
rect 14403 6554 14418 6754
rect 14970 6554 14985 6754
rect 15014 6554 15029 6754
rect 15581 6554 15596 6754
rect 15625 6554 15640 6754
rect 12559 5904 12574 6104
rect 12603 5904 12618 6104
rect 13170 5904 13185 6104
rect 13214 5904 13229 6104
rect 13781 5904 13796 6104
rect 13825 5904 13840 6104
rect 14359 5904 14374 6104
rect 14403 5904 14418 6104
rect 14970 5904 14985 6104
rect 15014 5904 15029 6104
rect 15581 5904 15596 6104
rect 15625 5904 15640 6104
rect 12559 5254 12574 5454
rect 12603 5254 12618 5454
rect 13170 5254 13185 5454
rect 13214 5254 13229 5454
rect 13781 5254 13796 5454
rect 13825 5254 13840 5454
rect 14359 5254 14374 5454
rect 14403 5254 14418 5454
rect 14970 5254 14985 5454
rect 15014 5254 15029 5454
rect 15581 5254 15596 5454
rect 15625 5254 15640 5454
rect 12559 4614 12574 4814
rect 12603 4614 12618 4814
rect 13170 4614 13185 4814
rect 13214 4614 13229 4814
rect 13781 4614 13796 4814
rect 13825 4614 13840 4814
rect 14359 4614 14374 4814
rect 14403 4614 14418 4814
rect 14970 4614 14985 4814
rect 15014 4614 15029 4814
rect 15581 4614 15596 4814
rect 15625 4614 15640 4814
<< ndiff >>
rect 13061 7663 13090 7670
rect 13061 7646 13067 7663
rect 13084 7646 13090 7663
rect 13061 7629 13090 7646
rect 13061 7612 13067 7629
rect 13084 7612 13090 7629
rect 13061 7595 13090 7612
rect 13061 7578 13067 7595
rect 13084 7578 13090 7595
rect 13061 7570 13090 7578
rect 13105 7570 13126 7670
rect 13141 7663 13170 7670
rect 13141 7646 13147 7663
rect 13164 7646 13170 7663
rect 13141 7629 13170 7646
rect 13141 7612 13147 7629
rect 13164 7612 13170 7629
rect 13141 7595 13170 7612
rect 13141 7578 13147 7595
rect 13164 7578 13170 7595
rect 13141 7570 13170 7578
rect 13185 7663 13214 7670
rect 13185 7646 13191 7663
rect 13208 7646 13214 7663
rect 13185 7629 13214 7646
rect 13185 7612 13191 7629
rect 13208 7612 13214 7629
rect 13185 7595 13214 7612
rect 13185 7578 13191 7595
rect 13208 7578 13214 7595
rect 13185 7570 13214 7578
rect 13229 7663 13258 7670
rect 13229 7646 13235 7663
rect 13252 7646 13258 7663
rect 13229 7629 13258 7646
rect 13229 7612 13235 7629
rect 13252 7612 13258 7629
rect 13229 7595 13258 7612
rect 13229 7578 13235 7595
rect 13252 7578 13258 7595
rect 13229 7570 13258 7578
rect 13273 7570 13294 7670
rect 13309 7663 13338 7670
rect 13309 7646 13315 7663
rect 13332 7646 13338 7663
rect 13309 7629 13338 7646
rect 13309 7612 13315 7629
rect 13332 7612 13338 7629
rect 13309 7595 13338 7612
rect 13309 7578 13315 7595
rect 13332 7578 13338 7595
rect 13309 7570 13338 7578
rect 13672 7663 13701 7670
rect 13672 7646 13678 7663
rect 13695 7646 13701 7663
rect 13672 7629 13701 7646
rect 13672 7612 13678 7629
rect 13695 7612 13701 7629
rect 13672 7595 13701 7612
rect 13672 7578 13678 7595
rect 13695 7578 13701 7595
rect 13672 7570 13701 7578
rect 13716 7570 13737 7670
rect 13752 7663 13781 7670
rect 13752 7646 13758 7663
rect 13775 7646 13781 7663
rect 13752 7629 13781 7646
rect 13752 7612 13758 7629
rect 13775 7612 13781 7629
rect 13752 7595 13781 7612
rect 13752 7578 13758 7595
rect 13775 7578 13781 7595
rect 13752 7570 13781 7578
rect 13796 7663 13825 7670
rect 13796 7646 13802 7663
rect 13819 7646 13825 7663
rect 13796 7629 13825 7646
rect 13796 7612 13802 7629
rect 13819 7612 13825 7629
rect 13796 7595 13825 7612
rect 13796 7578 13802 7595
rect 13819 7578 13825 7595
rect 13796 7570 13825 7578
rect 13840 7663 13869 7670
rect 13840 7646 13846 7663
rect 13863 7646 13869 7663
rect 13840 7629 13869 7646
rect 13840 7612 13846 7629
rect 13863 7612 13869 7629
rect 13840 7595 13869 7612
rect 13840 7578 13846 7595
rect 13863 7578 13869 7595
rect 13840 7570 13869 7578
rect 13884 7570 13905 7670
rect 13920 7663 13949 7670
rect 13920 7646 13926 7663
rect 13943 7646 13949 7663
rect 13920 7629 13949 7646
rect 13920 7612 13926 7629
rect 13943 7612 13949 7629
rect 13920 7595 13949 7612
rect 13920 7578 13926 7595
rect 13943 7578 13949 7595
rect 13920 7570 13949 7578
rect 14250 7663 14279 7670
rect 14250 7646 14256 7663
rect 14273 7646 14279 7663
rect 14250 7629 14279 7646
rect 14250 7612 14256 7629
rect 14273 7612 14279 7629
rect 14250 7595 14279 7612
rect 14250 7578 14256 7595
rect 14273 7578 14279 7595
rect 14250 7570 14279 7578
rect 14294 7570 14315 7670
rect 14330 7663 14359 7670
rect 14330 7646 14336 7663
rect 14353 7646 14359 7663
rect 14330 7629 14359 7646
rect 14330 7612 14336 7629
rect 14353 7612 14359 7629
rect 14330 7595 14359 7612
rect 14330 7578 14336 7595
rect 14353 7578 14359 7595
rect 14330 7570 14359 7578
rect 14374 7663 14403 7670
rect 14374 7646 14380 7663
rect 14397 7646 14403 7663
rect 14374 7629 14403 7646
rect 14374 7612 14380 7629
rect 14397 7612 14403 7629
rect 14374 7595 14403 7612
rect 14374 7578 14380 7595
rect 14397 7578 14403 7595
rect 14374 7570 14403 7578
rect 14418 7663 14447 7670
rect 14418 7646 14424 7663
rect 14441 7646 14447 7663
rect 14418 7629 14447 7646
rect 14418 7612 14424 7629
rect 14441 7612 14447 7629
rect 14418 7595 14447 7612
rect 14418 7578 14424 7595
rect 14441 7578 14447 7595
rect 14418 7570 14447 7578
rect 14462 7570 14483 7670
rect 14498 7663 14527 7670
rect 14498 7646 14504 7663
rect 14521 7646 14527 7663
rect 14498 7629 14527 7646
rect 14498 7612 14504 7629
rect 14521 7612 14527 7629
rect 14498 7595 14527 7612
rect 14498 7578 14504 7595
rect 14521 7578 14527 7595
rect 14498 7570 14527 7578
rect 14861 7663 14890 7670
rect 14861 7646 14867 7663
rect 14884 7646 14890 7663
rect 14861 7629 14890 7646
rect 14861 7612 14867 7629
rect 14884 7612 14890 7629
rect 14861 7595 14890 7612
rect 14861 7578 14867 7595
rect 14884 7578 14890 7595
rect 14861 7570 14890 7578
rect 14905 7570 14926 7670
rect 14941 7663 14970 7670
rect 14941 7646 14947 7663
rect 14964 7646 14970 7663
rect 14941 7629 14970 7646
rect 14941 7612 14947 7629
rect 14964 7612 14970 7629
rect 14941 7595 14970 7612
rect 14941 7578 14947 7595
rect 14964 7578 14970 7595
rect 14941 7570 14970 7578
rect 14985 7663 15014 7670
rect 14985 7646 14991 7663
rect 15008 7646 15014 7663
rect 14985 7629 15014 7646
rect 14985 7612 14991 7629
rect 15008 7612 15014 7629
rect 14985 7595 15014 7612
rect 14985 7578 14991 7595
rect 15008 7578 15014 7595
rect 14985 7570 15014 7578
rect 15029 7663 15058 7670
rect 15029 7646 15035 7663
rect 15052 7646 15058 7663
rect 15029 7629 15058 7646
rect 15029 7612 15035 7629
rect 15052 7612 15058 7629
rect 15029 7595 15058 7612
rect 15029 7578 15035 7595
rect 15052 7578 15058 7595
rect 15029 7570 15058 7578
rect 15073 7570 15094 7670
rect 15109 7663 15138 7670
rect 15109 7646 15115 7663
rect 15132 7646 15138 7663
rect 15109 7629 15138 7646
rect 15109 7612 15115 7629
rect 15132 7612 15138 7629
rect 15109 7595 15138 7612
rect 15109 7578 15115 7595
rect 15132 7578 15138 7595
rect 15109 7570 15138 7578
rect 15472 7663 15501 7670
rect 15472 7646 15478 7663
rect 15495 7646 15501 7663
rect 15472 7629 15501 7646
rect 15472 7612 15478 7629
rect 15495 7612 15501 7629
rect 15472 7595 15501 7612
rect 15472 7578 15478 7595
rect 15495 7578 15501 7595
rect 15472 7570 15501 7578
rect 15516 7570 15537 7670
rect 15552 7663 15581 7670
rect 15552 7646 15558 7663
rect 15575 7646 15581 7663
rect 15552 7629 15581 7646
rect 15552 7612 15558 7629
rect 15575 7612 15581 7629
rect 15552 7595 15581 7612
rect 15552 7578 15558 7595
rect 15575 7578 15581 7595
rect 15552 7570 15581 7578
rect 15596 7663 15625 7670
rect 15596 7646 15602 7663
rect 15619 7646 15625 7663
rect 15596 7629 15625 7646
rect 15596 7612 15602 7629
rect 15619 7612 15625 7629
rect 15596 7595 15625 7612
rect 15596 7578 15602 7595
rect 15619 7578 15625 7595
rect 15596 7570 15625 7578
rect 15640 7663 15669 7670
rect 15640 7646 15646 7663
rect 15663 7646 15669 7663
rect 15640 7629 15669 7646
rect 15640 7612 15646 7629
rect 15663 7612 15669 7629
rect 15640 7595 15669 7612
rect 15640 7578 15646 7595
rect 15663 7578 15669 7595
rect 15640 7570 15669 7578
rect 15684 7570 15705 7670
rect 15720 7663 15749 7670
rect 15720 7646 15726 7663
rect 15743 7646 15749 7663
rect 15720 7629 15749 7646
rect 15720 7612 15726 7629
rect 15743 7612 15749 7629
rect 15720 7595 15749 7612
rect 15720 7578 15726 7595
rect 15743 7578 15749 7595
rect 15720 7570 15749 7578
rect 12450 7013 12479 7020
rect 12450 6996 12456 7013
rect 12473 6996 12479 7013
rect 12450 6979 12479 6996
rect 12450 6962 12456 6979
rect 12473 6962 12479 6979
rect 12450 6945 12479 6962
rect 12450 6928 12456 6945
rect 12473 6928 12479 6945
rect 12450 6920 12479 6928
rect 12494 6920 12515 7020
rect 12530 7013 12559 7020
rect 12530 6996 12536 7013
rect 12553 6996 12559 7013
rect 12530 6979 12559 6996
rect 12530 6962 12536 6979
rect 12553 6962 12559 6979
rect 12530 6945 12559 6962
rect 12530 6928 12536 6945
rect 12553 6928 12559 6945
rect 12530 6920 12559 6928
rect 12574 7013 12603 7020
rect 12574 6996 12580 7013
rect 12597 6996 12603 7013
rect 12574 6979 12603 6996
rect 12574 6962 12580 6979
rect 12597 6962 12603 6979
rect 12574 6945 12603 6962
rect 12574 6928 12580 6945
rect 12597 6928 12603 6945
rect 12574 6920 12603 6928
rect 12618 7013 12647 7020
rect 12618 6996 12624 7013
rect 12641 6996 12647 7013
rect 12618 6979 12647 6996
rect 12618 6962 12624 6979
rect 12641 6962 12647 6979
rect 12618 6945 12647 6962
rect 12618 6928 12624 6945
rect 12641 6928 12647 6945
rect 12618 6920 12647 6928
rect 12662 6920 12683 7020
rect 12698 7013 12727 7020
rect 12698 6996 12704 7013
rect 12721 6996 12727 7013
rect 12698 6979 12727 6996
rect 12698 6962 12704 6979
rect 12721 6962 12727 6979
rect 12698 6945 12727 6962
rect 12698 6928 12704 6945
rect 12721 6928 12727 6945
rect 12698 6920 12727 6928
rect 13061 7013 13090 7020
rect 13061 6996 13067 7013
rect 13084 6996 13090 7013
rect 13061 6979 13090 6996
rect 13061 6962 13067 6979
rect 13084 6962 13090 6979
rect 13061 6945 13090 6962
rect 13061 6928 13067 6945
rect 13084 6928 13090 6945
rect 13061 6920 13090 6928
rect 13105 6920 13126 7020
rect 13141 7013 13170 7020
rect 13141 6996 13147 7013
rect 13164 6996 13170 7013
rect 13141 6979 13170 6996
rect 13141 6962 13147 6979
rect 13164 6962 13170 6979
rect 13141 6945 13170 6962
rect 13141 6928 13147 6945
rect 13164 6928 13170 6945
rect 13141 6920 13170 6928
rect 13185 7013 13214 7020
rect 13185 6996 13191 7013
rect 13208 6996 13214 7013
rect 13185 6979 13214 6996
rect 13185 6962 13191 6979
rect 13208 6962 13214 6979
rect 13185 6945 13214 6962
rect 13185 6928 13191 6945
rect 13208 6928 13214 6945
rect 13185 6920 13214 6928
rect 13229 7013 13258 7020
rect 13229 6996 13235 7013
rect 13252 6996 13258 7013
rect 13229 6979 13258 6996
rect 13229 6962 13235 6979
rect 13252 6962 13258 6979
rect 13229 6945 13258 6962
rect 13229 6928 13235 6945
rect 13252 6928 13258 6945
rect 13229 6920 13258 6928
rect 13273 6920 13294 7020
rect 13309 7013 13338 7020
rect 13309 6996 13315 7013
rect 13332 6996 13338 7013
rect 13309 6979 13338 6996
rect 13309 6962 13315 6979
rect 13332 6962 13338 6979
rect 13309 6945 13338 6962
rect 13309 6928 13315 6945
rect 13332 6928 13338 6945
rect 13309 6920 13338 6928
rect 13672 7013 13701 7020
rect 13672 6996 13678 7013
rect 13695 6996 13701 7013
rect 13672 6979 13701 6996
rect 13672 6962 13678 6979
rect 13695 6962 13701 6979
rect 13672 6945 13701 6962
rect 13672 6928 13678 6945
rect 13695 6928 13701 6945
rect 13672 6920 13701 6928
rect 13716 6920 13737 7020
rect 13752 7013 13781 7020
rect 13752 6996 13758 7013
rect 13775 6996 13781 7013
rect 13752 6979 13781 6996
rect 13752 6962 13758 6979
rect 13775 6962 13781 6979
rect 13752 6945 13781 6962
rect 13752 6928 13758 6945
rect 13775 6928 13781 6945
rect 13752 6920 13781 6928
rect 13796 7013 13825 7020
rect 13796 6996 13802 7013
rect 13819 6996 13825 7013
rect 13796 6979 13825 6996
rect 13796 6962 13802 6979
rect 13819 6962 13825 6979
rect 13796 6945 13825 6962
rect 13796 6928 13802 6945
rect 13819 6928 13825 6945
rect 13796 6920 13825 6928
rect 13840 7013 13869 7020
rect 13840 6996 13846 7013
rect 13863 6996 13869 7013
rect 13840 6979 13869 6996
rect 13840 6962 13846 6979
rect 13863 6962 13869 6979
rect 13840 6945 13869 6962
rect 13840 6928 13846 6945
rect 13863 6928 13869 6945
rect 13840 6920 13869 6928
rect 13884 6920 13905 7020
rect 13920 7013 13949 7020
rect 13920 6996 13926 7013
rect 13943 6996 13949 7013
rect 13920 6979 13949 6996
rect 13920 6962 13926 6979
rect 13943 6962 13949 6979
rect 13920 6945 13949 6962
rect 13920 6928 13926 6945
rect 13943 6928 13949 6945
rect 13920 6920 13949 6928
rect 14250 7013 14279 7020
rect 14250 6996 14256 7013
rect 14273 6996 14279 7013
rect 14250 6979 14279 6996
rect 14250 6962 14256 6979
rect 14273 6962 14279 6979
rect 14250 6945 14279 6962
rect 14250 6928 14256 6945
rect 14273 6928 14279 6945
rect 14250 6920 14279 6928
rect 14294 6920 14315 7020
rect 14330 7013 14359 7020
rect 14330 6996 14336 7013
rect 14353 6996 14359 7013
rect 14330 6979 14359 6996
rect 14330 6962 14336 6979
rect 14353 6962 14359 6979
rect 14330 6945 14359 6962
rect 14330 6928 14336 6945
rect 14353 6928 14359 6945
rect 14330 6920 14359 6928
rect 14374 7013 14403 7020
rect 14374 6996 14380 7013
rect 14397 6996 14403 7013
rect 14374 6979 14403 6996
rect 14374 6962 14380 6979
rect 14397 6962 14403 6979
rect 14374 6945 14403 6962
rect 14374 6928 14380 6945
rect 14397 6928 14403 6945
rect 14374 6920 14403 6928
rect 14418 7013 14447 7020
rect 14418 6996 14424 7013
rect 14441 6996 14447 7013
rect 14418 6979 14447 6996
rect 14418 6962 14424 6979
rect 14441 6962 14447 6979
rect 14418 6945 14447 6962
rect 14418 6928 14424 6945
rect 14441 6928 14447 6945
rect 14418 6920 14447 6928
rect 14462 6920 14483 7020
rect 14498 7013 14527 7020
rect 14498 6996 14504 7013
rect 14521 6996 14527 7013
rect 14498 6979 14527 6996
rect 14498 6962 14504 6979
rect 14521 6962 14527 6979
rect 14498 6945 14527 6962
rect 14498 6928 14504 6945
rect 14521 6928 14527 6945
rect 14498 6920 14527 6928
rect 14861 7013 14890 7020
rect 14861 6996 14867 7013
rect 14884 6996 14890 7013
rect 14861 6979 14890 6996
rect 14861 6962 14867 6979
rect 14884 6962 14890 6979
rect 14861 6945 14890 6962
rect 14861 6928 14867 6945
rect 14884 6928 14890 6945
rect 14861 6920 14890 6928
rect 14905 6920 14926 7020
rect 14941 7013 14970 7020
rect 14941 6996 14947 7013
rect 14964 6996 14970 7013
rect 14941 6979 14970 6996
rect 14941 6962 14947 6979
rect 14964 6962 14970 6979
rect 14941 6945 14970 6962
rect 14941 6928 14947 6945
rect 14964 6928 14970 6945
rect 14941 6920 14970 6928
rect 14985 7013 15014 7020
rect 14985 6996 14991 7013
rect 15008 6996 15014 7013
rect 14985 6979 15014 6996
rect 14985 6962 14991 6979
rect 15008 6962 15014 6979
rect 14985 6945 15014 6962
rect 14985 6928 14991 6945
rect 15008 6928 15014 6945
rect 14985 6920 15014 6928
rect 15029 7013 15058 7020
rect 15029 6996 15035 7013
rect 15052 6996 15058 7013
rect 15029 6979 15058 6996
rect 15029 6962 15035 6979
rect 15052 6962 15058 6979
rect 15029 6945 15058 6962
rect 15029 6928 15035 6945
rect 15052 6928 15058 6945
rect 15029 6920 15058 6928
rect 15073 6920 15094 7020
rect 15109 7013 15138 7020
rect 15109 6996 15115 7013
rect 15132 6996 15138 7013
rect 15109 6979 15138 6996
rect 15109 6962 15115 6979
rect 15132 6962 15138 6979
rect 15109 6945 15138 6962
rect 15109 6928 15115 6945
rect 15132 6928 15138 6945
rect 15109 6920 15138 6928
rect 15472 7013 15501 7020
rect 15472 6996 15478 7013
rect 15495 6996 15501 7013
rect 15472 6979 15501 6996
rect 15472 6962 15478 6979
rect 15495 6962 15501 6979
rect 15472 6945 15501 6962
rect 15472 6928 15478 6945
rect 15495 6928 15501 6945
rect 15472 6920 15501 6928
rect 15516 6920 15537 7020
rect 15552 7013 15581 7020
rect 15552 6996 15558 7013
rect 15575 6996 15581 7013
rect 15552 6979 15581 6996
rect 15552 6962 15558 6979
rect 15575 6962 15581 6979
rect 15552 6945 15581 6962
rect 15552 6928 15558 6945
rect 15575 6928 15581 6945
rect 15552 6920 15581 6928
rect 15596 7013 15625 7020
rect 15596 6996 15602 7013
rect 15619 6996 15625 7013
rect 15596 6979 15625 6996
rect 15596 6962 15602 6979
rect 15619 6962 15625 6979
rect 15596 6945 15625 6962
rect 15596 6928 15602 6945
rect 15619 6928 15625 6945
rect 15596 6920 15625 6928
rect 15640 7013 15669 7020
rect 15640 6996 15646 7013
rect 15663 6996 15669 7013
rect 15640 6979 15669 6996
rect 15640 6962 15646 6979
rect 15663 6962 15669 6979
rect 15640 6945 15669 6962
rect 15640 6928 15646 6945
rect 15663 6928 15669 6945
rect 15640 6920 15669 6928
rect 15684 6920 15705 7020
rect 15720 7013 15749 7020
rect 15720 6996 15726 7013
rect 15743 6996 15749 7013
rect 15720 6979 15749 6996
rect 15720 6962 15726 6979
rect 15743 6962 15749 6979
rect 15720 6945 15749 6962
rect 15720 6928 15726 6945
rect 15743 6928 15749 6945
rect 15720 6920 15749 6928
rect 12450 6373 12479 6380
rect 12450 6356 12456 6373
rect 12473 6356 12479 6373
rect 12450 6339 12479 6356
rect 12450 6322 12456 6339
rect 12473 6322 12479 6339
rect 12450 6305 12479 6322
rect 12450 6288 12456 6305
rect 12473 6288 12479 6305
rect 12450 6280 12479 6288
rect 12494 6280 12515 6380
rect 12530 6373 12559 6380
rect 12530 6356 12536 6373
rect 12553 6356 12559 6373
rect 12530 6339 12559 6356
rect 12530 6322 12536 6339
rect 12553 6322 12559 6339
rect 12530 6305 12559 6322
rect 12530 6288 12536 6305
rect 12553 6288 12559 6305
rect 12530 6280 12559 6288
rect 12574 6373 12603 6380
rect 12574 6356 12580 6373
rect 12597 6356 12603 6373
rect 12574 6339 12603 6356
rect 12574 6322 12580 6339
rect 12597 6322 12603 6339
rect 12574 6305 12603 6322
rect 12574 6288 12580 6305
rect 12597 6288 12603 6305
rect 12574 6280 12603 6288
rect 12618 6373 12647 6380
rect 12618 6356 12624 6373
rect 12641 6356 12647 6373
rect 12618 6339 12647 6356
rect 12618 6322 12624 6339
rect 12641 6322 12647 6339
rect 12618 6305 12647 6322
rect 12618 6288 12624 6305
rect 12641 6288 12647 6305
rect 12618 6280 12647 6288
rect 12662 6280 12683 6380
rect 12698 6373 12727 6380
rect 12698 6356 12704 6373
rect 12721 6356 12727 6373
rect 12698 6339 12727 6356
rect 12698 6322 12704 6339
rect 12721 6322 12727 6339
rect 12698 6305 12727 6322
rect 12698 6288 12704 6305
rect 12721 6288 12727 6305
rect 12698 6280 12727 6288
rect 13061 6373 13090 6380
rect 13061 6356 13067 6373
rect 13084 6356 13090 6373
rect 13061 6339 13090 6356
rect 13061 6322 13067 6339
rect 13084 6322 13090 6339
rect 13061 6305 13090 6322
rect 13061 6288 13067 6305
rect 13084 6288 13090 6305
rect 13061 6280 13090 6288
rect 13105 6280 13126 6380
rect 13141 6373 13170 6380
rect 13141 6356 13147 6373
rect 13164 6356 13170 6373
rect 13141 6339 13170 6356
rect 13141 6322 13147 6339
rect 13164 6322 13170 6339
rect 13141 6305 13170 6322
rect 13141 6288 13147 6305
rect 13164 6288 13170 6305
rect 13141 6280 13170 6288
rect 13185 6373 13214 6380
rect 13185 6356 13191 6373
rect 13208 6356 13214 6373
rect 13185 6339 13214 6356
rect 13185 6322 13191 6339
rect 13208 6322 13214 6339
rect 13185 6305 13214 6322
rect 13185 6288 13191 6305
rect 13208 6288 13214 6305
rect 13185 6280 13214 6288
rect 13229 6373 13258 6380
rect 13229 6356 13235 6373
rect 13252 6356 13258 6373
rect 13229 6339 13258 6356
rect 13229 6322 13235 6339
rect 13252 6322 13258 6339
rect 13229 6305 13258 6322
rect 13229 6288 13235 6305
rect 13252 6288 13258 6305
rect 13229 6280 13258 6288
rect 13273 6280 13294 6380
rect 13309 6373 13338 6380
rect 13309 6356 13315 6373
rect 13332 6356 13338 6373
rect 13309 6339 13338 6356
rect 13309 6322 13315 6339
rect 13332 6322 13338 6339
rect 13309 6305 13338 6322
rect 13309 6288 13315 6305
rect 13332 6288 13338 6305
rect 13309 6280 13338 6288
rect 13672 6373 13701 6380
rect 13672 6356 13678 6373
rect 13695 6356 13701 6373
rect 13672 6339 13701 6356
rect 13672 6322 13678 6339
rect 13695 6322 13701 6339
rect 13672 6305 13701 6322
rect 13672 6288 13678 6305
rect 13695 6288 13701 6305
rect 13672 6280 13701 6288
rect 13716 6280 13737 6380
rect 13752 6373 13781 6380
rect 13752 6356 13758 6373
rect 13775 6356 13781 6373
rect 13752 6339 13781 6356
rect 13752 6322 13758 6339
rect 13775 6322 13781 6339
rect 13752 6305 13781 6322
rect 13752 6288 13758 6305
rect 13775 6288 13781 6305
rect 13752 6280 13781 6288
rect 13796 6373 13825 6380
rect 13796 6356 13802 6373
rect 13819 6356 13825 6373
rect 13796 6339 13825 6356
rect 13796 6322 13802 6339
rect 13819 6322 13825 6339
rect 13796 6305 13825 6322
rect 13796 6288 13802 6305
rect 13819 6288 13825 6305
rect 13796 6280 13825 6288
rect 13840 6373 13869 6380
rect 13840 6356 13846 6373
rect 13863 6356 13869 6373
rect 13840 6339 13869 6356
rect 13840 6322 13846 6339
rect 13863 6322 13869 6339
rect 13840 6305 13869 6322
rect 13840 6288 13846 6305
rect 13863 6288 13869 6305
rect 13840 6280 13869 6288
rect 13884 6280 13905 6380
rect 13920 6373 13949 6380
rect 13920 6356 13926 6373
rect 13943 6356 13949 6373
rect 13920 6339 13949 6356
rect 13920 6322 13926 6339
rect 13943 6322 13949 6339
rect 13920 6305 13949 6322
rect 13920 6288 13926 6305
rect 13943 6288 13949 6305
rect 13920 6280 13949 6288
rect 14250 6373 14279 6380
rect 14250 6356 14256 6373
rect 14273 6356 14279 6373
rect 14250 6339 14279 6356
rect 14250 6322 14256 6339
rect 14273 6322 14279 6339
rect 14250 6305 14279 6322
rect 14250 6288 14256 6305
rect 14273 6288 14279 6305
rect 14250 6280 14279 6288
rect 14294 6280 14315 6380
rect 14330 6373 14359 6380
rect 14330 6356 14336 6373
rect 14353 6356 14359 6373
rect 14330 6339 14359 6356
rect 14330 6322 14336 6339
rect 14353 6322 14359 6339
rect 14330 6305 14359 6322
rect 14330 6288 14336 6305
rect 14353 6288 14359 6305
rect 14330 6280 14359 6288
rect 14374 6373 14403 6380
rect 14374 6356 14380 6373
rect 14397 6356 14403 6373
rect 14374 6339 14403 6356
rect 14374 6322 14380 6339
rect 14397 6322 14403 6339
rect 14374 6305 14403 6322
rect 14374 6288 14380 6305
rect 14397 6288 14403 6305
rect 14374 6280 14403 6288
rect 14418 6373 14447 6380
rect 14418 6356 14424 6373
rect 14441 6356 14447 6373
rect 14418 6339 14447 6356
rect 14418 6322 14424 6339
rect 14441 6322 14447 6339
rect 14418 6305 14447 6322
rect 14418 6288 14424 6305
rect 14441 6288 14447 6305
rect 14418 6280 14447 6288
rect 14462 6280 14483 6380
rect 14498 6373 14527 6380
rect 14498 6356 14504 6373
rect 14521 6356 14527 6373
rect 14498 6339 14527 6356
rect 14498 6322 14504 6339
rect 14521 6322 14527 6339
rect 14498 6305 14527 6322
rect 14498 6288 14504 6305
rect 14521 6288 14527 6305
rect 14498 6280 14527 6288
rect 14861 6373 14890 6380
rect 14861 6356 14867 6373
rect 14884 6356 14890 6373
rect 14861 6339 14890 6356
rect 14861 6322 14867 6339
rect 14884 6322 14890 6339
rect 14861 6305 14890 6322
rect 14861 6288 14867 6305
rect 14884 6288 14890 6305
rect 14861 6280 14890 6288
rect 14905 6280 14926 6380
rect 14941 6373 14970 6380
rect 14941 6356 14947 6373
rect 14964 6356 14970 6373
rect 14941 6339 14970 6356
rect 14941 6322 14947 6339
rect 14964 6322 14970 6339
rect 14941 6305 14970 6322
rect 14941 6288 14947 6305
rect 14964 6288 14970 6305
rect 14941 6280 14970 6288
rect 14985 6373 15014 6380
rect 14985 6356 14991 6373
rect 15008 6356 15014 6373
rect 14985 6339 15014 6356
rect 14985 6322 14991 6339
rect 15008 6322 15014 6339
rect 14985 6305 15014 6322
rect 14985 6288 14991 6305
rect 15008 6288 15014 6305
rect 14985 6280 15014 6288
rect 15029 6373 15058 6380
rect 15029 6356 15035 6373
rect 15052 6356 15058 6373
rect 15029 6339 15058 6356
rect 15029 6322 15035 6339
rect 15052 6322 15058 6339
rect 15029 6305 15058 6322
rect 15029 6288 15035 6305
rect 15052 6288 15058 6305
rect 15029 6280 15058 6288
rect 15073 6280 15094 6380
rect 15109 6373 15138 6380
rect 15109 6356 15115 6373
rect 15132 6356 15138 6373
rect 15109 6339 15138 6356
rect 15109 6322 15115 6339
rect 15132 6322 15138 6339
rect 15109 6305 15138 6322
rect 15109 6288 15115 6305
rect 15132 6288 15138 6305
rect 15109 6280 15138 6288
rect 15472 6373 15501 6380
rect 15472 6356 15478 6373
rect 15495 6356 15501 6373
rect 15472 6339 15501 6356
rect 15472 6322 15478 6339
rect 15495 6322 15501 6339
rect 15472 6305 15501 6322
rect 15472 6288 15478 6305
rect 15495 6288 15501 6305
rect 15472 6280 15501 6288
rect 15516 6280 15537 6380
rect 15552 6373 15581 6380
rect 15552 6356 15558 6373
rect 15575 6356 15581 6373
rect 15552 6339 15581 6356
rect 15552 6322 15558 6339
rect 15575 6322 15581 6339
rect 15552 6305 15581 6322
rect 15552 6288 15558 6305
rect 15575 6288 15581 6305
rect 15552 6280 15581 6288
rect 15596 6373 15625 6380
rect 15596 6356 15602 6373
rect 15619 6356 15625 6373
rect 15596 6339 15625 6356
rect 15596 6322 15602 6339
rect 15619 6322 15625 6339
rect 15596 6305 15625 6322
rect 15596 6288 15602 6305
rect 15619 6288 15625 6305
rect 15596 6280 15625 6288
rect 15640 6373 15669 6380
rect 15640 6356 15646 6373
rect 15663 6356 15669 6373
rect 15640 6339 15669 6356
rect 15640 6322 15646 6339
rect 15663 6322 15669 6339
rect 15640 6305 15669 6322
rect 15640 6288 15646 6305
rect 15663 6288 15669 6305
rect 15640 6280 15669 6288
rect 15684 6280 15705 6380
rect 15720 6373 15749 6380
rect 15720 6356 15726 6373
rect 15743 6356 15749 6373
rect 15720 6339 15749 6356
rect 15720 6322 15726 6339
rect 15743 6322 15749 6339
rect 15720 6305 15749 6322
rect 15720 6288 15726 6305
rect 15743 6288 15749 6305
rect 15720 6280 15749 6288
rect 12450 5723 12479 5730
rect 12450 5706 12456 5723
rect 12473 5706 12479 5723
rect 12450 5689 12479 5706
rect 12450 5672 12456 5689
rect 12473 5672 12479 5689
rect 12450 5655 12479 5672
rect 12450 5638 12456 5655
rect 12473 5638 12479 5655
rect 12450 5630 12479 5638
rect 12494 5630 12515 5730
rect 12530 5723 12559 5730
rect 12530 5706 12536 5723
rect 12553 5706 12559 5723
rect 12530 5689 12559 5706
rect 12530 5672 12536 5689
rect 12553 5672 12559 5689
rect 12530 5655 12559 5672
rect 12530 5638 12536 5655
rect 12553 5638 12559 5655
rect 12530 5630 12559 5638
rect 12574 5723 12603 5730
rect 12574 5706 12580 5723
rect 12597 5706 12603 5723
rect 12574 5689 12603 5706
rect 12574 5672 12580 5689
rect 12597 5672 12603 5689
rect 12574 5655 12603 5672
rect 12574 5638 12580 5655
rect 12597 5638 12603 5655
rect 12574 5630 12603 5638
rect 12618 5723 12647 5730
rect 12618 5706 12624 5723
rect 12641 5706 12647 5723
rect 12618 5689 12647 5706
rect 12618 5672 12624 5689
rect 12641 5672 12647 5689
rect 12618 5655 12647 5672
rect 12618 5638 12624 5655
rect 12641 5638 12647 5655
rect 12618 5630 12647 5638
rect 12662 5630 12683 5730
rect 12698 5723 12727 5730
rect 12698 5706 12704 5723
rect 12721 5706 12727 5723
rect 12698 5689 12727 5706
rect 12698 5672 12704 5689
rect 12721 5672 12727 5689
rect 12698 5655 12727 5672
rect 12698 5638 12704 5655
rect 12721 5638 12727 5655
rect 12698 5630 12727 5638
rect 13061 5723 13090 5730
rect 13061 5706 13067 5723
rect 13084 5706 13090 5723
rect 13061 5689 13090 5706
rect 13061 5672 13067 5689
rect 13084 5672 13090 5689
rect 13061 5655 13090 5672
rect 13061 5638 13067 5655
rect 13084 5638 13090 5655
rect 13061 5630 13090 5638
rect 13105 5630 13126 5730
rect 13141 5723 13170 5730
rect 13141 5706 13147 5723
rect 13164 5706 13170 5723
rect 13141 5689 13170 5706
rect 13141 5672 13147 5689
rect 13164 5672 13170 5689
rect 13141 5655 13170 5672
rect 13141 5638 13147 5655
rect 13164 5638 13170 5655
rect 13141 5630 13170 5638
rect 13185 5723 13214 5730
rect 13185 5706 13191 5723
rect 13208 5706 13214 5723
rect 13185 5689 13214 5706
rect 13185 5672 13191 5689
rect 13208 5672 13214 5689
rect 13185 5655 13214 5672
rect 13185 5638 13191 5655
rect 13208 5638 13214 5655
rect 13185 5630 13214 5638
rect 13229 5723 13258 5730
rect 13229 5706 13235 5723
rect 13252 5706 13258 5723
rect 13229 5689 13258 5706
rect 13229 5672 13235 5689
rect 13252 5672 13258 5689
rect 13229 5655 13258 5672
rect 13229 5638 13235 5655
rect 13252 5638 13258 5655
rect 13229 5630 13258 5638
rect 13273 5630 13294 5730
rect 13309 5723 13338 5730
rect 13309 5706 13315 5723
rect 13332 5706 13338 5723
rect 13309 5689 13338 5706
rect 13309 5672 13315 5689
rect 13332 5672 13338 5689
rect 13309 5655 13338 5672
rect 13309 5638 13315 5655
rect 13332 5638 13338 5655
rect 13309 5630 13338 5638
rect 13672 5723 13701 5730
rect 13672 5706 13678 5723
rect 13695 5706 13701 5723
rect 13672 5689 13701 5706
rect 13672 5672 13678 5689
rect 13695 5672 13701 5689
rect 13672 5655 13701 5672
rect 13672 5638 13678 5655
rect 13695 5638 13701 5655
rect 13672 5630 13701 5638
rect 13716 5630 13737 5730
rect 13752 5723 13781 5730
rect 13752 5706 13758 5723
rect 13775 5706 13781 5723
rect 13752 5689 13781 5706
rect 13752 5672 13758 5689
rect 13775 5672 13781 5689
rect 13752 5655 13781 5672
rect 13752 5638 13758 5655
rect 13775 5638 13781 5655
rect 13752 5630 13781 5638
rect 13796 5723 13825 5730
rect 13796 5706 13802 5723
rect 13819 5706 13825 5723
rect 13796 5689 13825 5706
rect 13796 5672 13802 5689
rect 13819 5672 13825 5689
rect 13796 5655 13825 5672
rect 13796 5638 13802 5655
rect 13819 5638 13825 5655
rect 13796 5630 13825 5638
rect 13840 5723 13869 5730
rect 13840 5706 13846 5723
rect 13863 5706 13869 5723
rect 13840 5689 13869 5706
rect 13840 5672 13846 5689
rect 13863 5672 13869 5689
rect 13840 5655 13869 5672
rect 13840 5638 13846 5655
rect 13863 5638 13869 5655
rect 13840 5630 13869 5638
rect 13884 5630 13905 5730
rect 13920 5723 13949 5730
rect 13920 5706 13926 5723
rect 13943 5706 13949 5723
rect 13920 5689 13949 5706
rect 13920 5672 13926 5689
rect 13943 5672 13949 5689
rect 13920 5655 13949 5672
rect 13920 5638 13926 5655
rect 13943 5638 13949 5655
rect 13920 5630 13949 5638
rect 14250 5723 14279 5730
rect 14250 5706 14256 5723
rect 14273 5706 14279 5723
rect 14250 5689 14279 5706
rect 14250 5672 14256 5689
rect 14273 5672 14279 5689
rect 14250 5655 14279 5672
rect 14250 5638 14256 5655
rect 14273 5638 14279 5655
rect 14250 5630 14279 5638
rect 14294 5630 14315 5730
rect 14330 5723 14359 5730
rect 14330 5706 14336 5723
rect 14353 5706 14359 5723
rect 14330 5689 14359 5706
rect 14330 5672 14336 5689
rect 14353 5672 14359 5689
rect 14330 5655 14359 5672
rect 14330 5638 14336 5655
rect 14353 5638 14359 5655
rect 14330 5630 14359 5638
rect 14374 5723 14403 5730
rect 14374 5706 14380 5723
rect 14397 5706 14403 5723
rect 14374 5689 14403 5706
rect 14374 5672 14380 5689
rect 14397 5672 14403 5689
rect 14374 5655 14403 5672
rect 14374 5638 14380 5655
rect 14397 5638 14403 5655
rect 14374 5630 14403 5638
rect 14418 5723 14447 5730
rect 14418 5706 14424 5723
rect 14441 5706 14447 5723
rect 14418 5689 14447 5706
rect 14418 5672 14424 5689
rect 14441 5672 14447 5689
rect 14418 5655 14447 5672
rect 14418 5638 14424 5655
rect 14441 5638 14447 5655
rect 14418 5630 14447 5638
rect 14462 5630 14483 5730
rect 14498 5723 14527 5730
rect 14498 5706 14504 5723
rect 14521 5706 14527 5723
rect 14498 5689 14527 5706
rect 14498 5672 14504 5689
rect 14521 5672 14527 5689
rect 14498 5655 14527 5672
rect 14498 5638 14504 5655
rect 14521 5638 14527 5655
rect 14498 5630 14527 5638
rect 14861 5723 14890 5730
rect 14861 5706 14867 5723
rect 14884 5706 14890 5723
rect 14861 5689 14890 5706
rect 14861 5672 14867 5689
rect 14884 5672 14890 5689
rect 14861 5655 14890 5672
rect 14861 5638 14867 5655
rect 14884 5638 14890 5655
rect 14861 5630 14890 5638
rect 14905 5630 14926 5730
rect 14941 5723 14970 5730
rect 14941 5706 14947 5723
rect 14964 5706 14970 5723
rect 14941 5689 14970 5706
rect 14941 5672 14947 5689
rect 14964 5672 14970 5689
rect 14941 5655 14970 5672
rect 14941 5638 14947 5655
rect 14964 5638 14970 5655
rect 14941 5630 14970 5638
rect 14985 5723 15014 5730
rect 14985 5706 14991 5723
rect 15008 5706 15014 5723
rect 14985 5689 15014 5706
rect 14985 5672 14991 5689
rect 15008 5672 15014 5689
rect 14985 5655 15014 5672
rect 14985 5638 14991 5655
rect 15008 5638 15014 5655
rect 14985 5630 15014 5638
rect 15029 5723 15058 5730
rect 15029 5706 15035 5723
rect 15052 5706 15058 5723
rect 15029 5689 15058 5706
rect 15029 5672 15035 5689
rect 15052 5672 15058 5689
rect 15029 5655 15058 5672
rect 15029 5638 15035 5655
rect 15052 5638 15058 5655
rect 15029 5630 15058 5638
rect 15073 5630 15094 5730
rect 15109 5723 15138 5730
rect 15109 5706 15115 5723
rect 15132 5706 15138 5723
rect 15109 5689 15138 5706
rect 15109 5672 15115 5689
rect 15132 5672 15138 5689
rect 15109 5655 15138 5672
rect 15109 5638 15115 5655
rect 15132 5638 15138 5655
rect 15109 5630 15138 5638
rect 15472 5723 15501 5730
rect 15472 5706 15478 5723
rect 15495 5706 15501 5723
rect 15472 5689 15501 5706
rect 15472 5672 15478 5689
rect 15495 5672 15501 5689
rect 15472 5655 15501 5672
rect 15472 5638 15478 5655
rect 15495 5638 15501 5655
rect 15472 5630 15501 5638
rect 15516 5630 15537 5730
rect 15552 5723 15581 5730
rect 15552 5706 15558 5723
rect 15575 5706 15581 5723
rect 15552 5689 15581 5706
rect 15552 5672 15558 5689
rect 15575 5672 15581 5689
rect 15552 5655 15581 5672
rect 15552 5638 15558 5655
rect 15575 5638 15581 5655
rect 15552 5630 15581 5638
rect 15596 5723 15625 5730
rect 15596 5706 15602 5723
rect 15619 5706 15625 5723
rect 15596 5689 15625 5706
rect 15596 5672 15602 5689
rect 15619 5672 15625 5689
rect 15596 5655 15625 5672
rect 15596 5638 15602 5655
rect 15619 5638 15625 5655
rect 15596 5630 15625 5638
rect 15640 5723 15669 5730
rect 15640 5706 15646 5723
rect 15663 5706 15669 5723
rect 15640 5689 15669 5706
rect 15640 5672 15646 5689
rect 15663 5672 15669 5689
rect 15640 5655 15669 5672
rect 15640 5638 15646 5655
rect 15663 5638 15669 5655
rect 15640 5630 15669 5638
rect 15684 5630 15705 5730
rect 15720 5723 15749 5730
rect 15720 5706 15726 5723
rect 15743 5706 15749 5723
rect 15720 5689 15749 5706
rect 15720 5672 15726 5689
rect 15743 5672 15749 5689
rect 15720 5655 15749 5672
rect 15720 5638 15726 5655
rect 15743 5638 15749 5655
rect 15720 5630 15749 5638
rect 12450 5073 12479 5080
rect 12450 5056 12456 5073
rect 12473 5056 12479 5073
rect 12450 5039 12479 5056
rect 12450 5022 12456 5039
rect 12473 5022 12479 5039
rect 12450 5005 12479 5022
rect 12450 4988 12456 5005
rect 12473 4988 12479 5005
rect 12450 4980 12479 4988
rect 12494 4980 12515 5080
rect 12530 5073 12559 5080
rect 12530 5056 12536 5073
rect 12553 5056 12559 5073
rect 12530 5039 12559 5056
rect 12530 5022 12536 5039
rect 12553 5022 12559 5039
rect 12530 5005 12559 5022
rect 12530 4988 12536 5005
rect 12553 4988 12559 5005
rect 12530 4980 12559 4988
rect 12574 5073 12603 5080
rect 12574 5056 12580 5073
rect 12597 5056 12603 5073
rect 12574 5039 12603 5056
rect 12574 5022 12580 5039
rect 12597 5022 12603 5039
rect 12574 5005 12603 5022
rect 12574 4988 12580 5005
rect 12597 4988 12603 5005
rect 12574 4980 12603 4988
rect 12618 5073 12647 5080
rect 12618 5056 12624 5073
rect 12641 5056 12647 5073
rect 12618 5039 12647 5056
rect 12618 5022 12624 5039
rect 12641 5022 12647 5039
rect 12618 5005 12647 5022
rect 12618 4988 12624 5005
rect 12641 4988 12647 5005
rect 12618 4980 12647 4988
rect 12662 4980 12683 5080
rect 12698 5073 12727 5080
rect 12698 5056 12704 5073
rect 12721 5056 12727 5073
rect 12698 5039 12727 5056
rect 12698 5022 12704 5039
rect 12721 5022 12727 5039
rect 12698 5005 12727 5022
rect 12698 4988 12704 5005
rect 12721 4988 12727 5005
rect 12698 4980 12727 4988
rect 13061 5073 13090 5080
rect 13061 5056 13067 5073
rect 13084 5056 13090 5073
rect 13061 5039 13090 5056
rect 13061 5022 13067 5039
rect 13084 5022 13090 5039
rect 13061 5005 13090 5022
rect 13061 4988 13067 5005
rect 13084 4988 13090 5005
rect 13061 4980 13090 4988
rect 13105 4980 13126 5080
rect 13141 5073 13170 5080
rect 13141 5056 13147 5073
rect 13164 5056 13170 5073
rect 13141 5039 13170 5056
rect 13141 5022 13147 5039
rect 13164 5022 13170 5039
rect 13141 5005 13170 5022
rect 13141 4988 13147 5005
rect 13164 4988 13170 5005
rect 13141 4980 13170 4988
rect 13185 5073 13214 5080
rect 13185 5056 13191 5073
rect 13208 5056 13214 5073
rect 13185 5039 13214 5056
rect 13185 5022 13191 5039
rect 13208 5022 13214 5039
rect 13185 5005 13214 5022
rect 13185 4988 13191 5005
rect 13208 4988 13214 5005
rect 13185 4980 13214 4988
rect 13229 5073 13258 5080
rect 13229 5056 13235 5073
rect 13252 5056 13258 5073
rect 13229 5039 13258 5056
rect 13229 5022 13235 5039
rect 13252 5022 13258 5039
rect 13229 5005 13258 5022
rect 13229 4988 13235 5005
rect 13252 4988 13258 5005
rect 13229 4980 13258 4988
rect 13273 4980 13294 5080
rect 13309 5073 13338 5080
rect 13309 5056 13315 5073
rect 13332 5056 13338 5073
rect 13309 5039 13338 5056
rect 13309 5022 13315 5039
rect 13332 5022 13338 5039
rect 13309 5005 13338 5022
rect 13309 4988 13315 5005
rect 13332 4988 13338 5005
rect 13309 4980 13338 4988
rect 13672 5073 13701 5080
rect 13672 5056 13678 5073
rect 13695 5056 13701 5073
rect 13672 5039 13701 5056
rect 13672 5022 13678 5039
rect 13695 5022 13701 5039
rect 13672 5005 13701 5022
rect 13672 4988 13678 5005
rect 13695 4988 13701 5005
rect 13672 4980 13701 4988
rect 13716 4980 13737 5080
rect 13752 5073 13781 5080
rect 13752 5056 13758 5073
rect 13775 5056 13781 5073
rect 13752 5039 13781 5056
rect 13752 5022 13758 5039
rect 13775 5022 13781 5039
rect 13752 5005 13781 5022
rect 13752 4988 13758 5005
rect 13775 4988 13781 5005
rect 13752 4980 13781 4988
rect 13796 5073 13825 5080
rect 13796 5056 13802 5073
rect 13819 5056 13825 5073
rect 13796 5039 13825 5056
rect 13796 5022 13802 5039
rect 13819 5022 13825 5039
rect 13796 5005 13825 5022
rect 13796 4988 13802 5005
rect 13819 4988 13825 5005
rect 13796 4980 13825 4988
rect 13840 5073 13869 5080
rect 13840 5056 13846 5073
rect 13863 5056 13869 5073
rect 13840 5039 13869 5056
rect 13840 5022 13846 5039
rect 13863 5022 13869 5039
rect 13840 5005 13869 5022
rect 13840 4988 13846 5005
rect 13863 4988 13869 5005
rect 13840 4980 13869 4988
rect 13884 4980 13905 5080
rect 13920 5073 13949 5080
rect 13920 5056 13926 5073
rect 13943 5056 13949 5073
rect 13920 5039 13949 5056
rect 13920 5022 13926 5039
rect 13943 5022 13949 5039
rect 13920 5005 13949 5022
rect 13920 4988 13926 5005
rect 13943 4988 13949 5005
rect 13920 4980 13949 4988
rect 14250 5073 14279 5080
rect 14250 5056 14256 5073
rect 14273 5056 14279 5073
rect 14250 5039 14279 5056
rect 14250 5022 14256 5039
rect 14273 5022 14279 5039
rect 14250 5005 14279 5022
rect 14250 4988 14256 5005
rect 14273 4988 14279 5005
rect 14250 4980 14279 4988
rect 14294 4980 14315 5080
rect 14330 5073 14359 5080
rect 14330 5056 14336 5073
rect 14353 5056 14359 5073
rect 14330 5039 14359 5056
rect 14330 5022 14336 5039
rect 14353 5022 14359 5039
rect 14330 5005 14359 5022
rect 14330 4988 14336 5005
rect 14353 4988 14359 5005
rect 14330 4980 14359 4988
rect 14374 5073 14403 5080
rect 14374 5056 14380 5073
rect 14397 5056 14403 5073
rect 14374 5039 14403 5056
rect 14374 5022 14380 5039
rect 14397 5022 14403 5039
rect 14374 5005 14403 5022
rect 14374 4988 14380 5005
rect 14397 4988 14403 5005
rect 14374 4980 14403 4988
rect 14418 5073 14447 5080
rect 14418 5056 14424 5073
rect 14441 5056 14447 5073
rect 14418 5039 14447 5056
rect 14418 5022 14424 5039
rect 14441 5022 14447 5039
rect 14418 5005 14447 5022
rect 14418 4988 14424 5005
rect 14441 4988 14447 5005
rect 14418 4980 14447 4988
rect 14462 4980 14483 5080
rect 14498 5073 14527 5080
rect 14498 5056 14504 5073
rect 14521 5056 14527 5073
rect 14498 5039 14527 5056
rect 14498 5022 14504 5039
rect 14521 5022 14527 5039
rect 14498 5005 14527 5022
rect 14498 4988 14504 5005
rect 14521 4988 14527 5005
rect 14498 4980 14527 4988
rect 14861 5073 14890 5080
rect 14861 5056 14867 5073
rect 14884 5056 14890 5073
rect 14861 5039 14890 5056
rect 14861 5022 14867 5039
rect 14884 5022 14890 5039
rect 14861 5005 14890 5022
rect 14861 4988 14867 5005
rect 14884 4988 14890 5005
rect 14861 4980 14890 4988
rect 14905 4980 14926 5080
rect 14941 5073 14970 5080
rect 14941 5056 14947 5073
rect 14964 5056 14970 5073
rect 14941 5039 14970 5056
rect 14941 5022 14947 5039
rect 14964 5022 14970 5039
rect 14941 5005 14970 5022
rect 14941 4988 14947 5005
rect 14964 4988 14970 5005
rect 14941 4980 14970 4988
rect 14985 5073 15014 5080
rect 14985 5056 14991 5073
rect 15008 5056 15014 5073
rect 14985 5039 15014 5056
rect 14985 5022 14991 5039
rect 15008 5022 15014 5039
rect 14985 5005 15014 5022
rect 14985 4988 14991 5005
rect 15008 4988 15014 5005
rect 14985 4980 15014 4988
rect 15029 5073 15058 5080
rect 15029 5056 15035 5073
rect 15052 5056 15058 5073
rect 15029 5039 15058 5056
rect 15029 5022 15035 5039
rect 15052 5022 15058 5039
rect 15029 5005 15058 5022
rect 15029 4988 15035 5005
rect 15052 4988 15058 5005
rect 15029 4980 15058 4988
rect 15073 4980 15094 5080
rect 15109 5073 15138 5080
rect 15109 5056 15115 5073
rect 15132 5056 15138 5073
rect 15109 5039 15138 5056
rect 15109 5022 15115 5039
rect 15132 5022 15138 5039
rect 15109 5005 15138 5022
rect 15109 4988 15115 5005
rect 15132 4988 15138 5005
rect 15109 4980 15138 4988
rect 15472 5073 15501 5080
rect 15472 5056 15478 5073
rect 15495 5056 15501 5073
rect 15472 5039 15501 5056
rect 15472 5022 15478 5039
rect 15495 5022 15501 5039
rect 15472 5005 15501 5022
rect 15472 4988 15478 5005
rect 15495 4988 15501 5005
rect 15472 4980 15501 4988
rect 15516 4980 15537 5080
rect 15552 5073 15581 5080
rect 15552 5056 15558 5073
rect 15575 5056 15581 5073
rect 15552 5039 15581 5056
rect 15552 5022 15558 5039
rect 15575 5022 15581 5039
rect 15552 5005 15581 5022
rect 15552 4988 15558 5005
rect 15575 4988 15581 5005
rect 15552 4980 15581 4988
rect 15596 5073 15625 5080
rect 15596 5056 15602 5073
rect 15619 5056 15625 5073
rect 15596 5039 15625 5056
rect 15596 5022 15602 5039
rect 15619 5022 15625 5039
rect 15596 5005 15625 5022
rect 15596 4988 15602 5005
rect 15619 4988 15625 5005
rect 15596 4980 15625 4988
rect 15640 5073 15669 5080
rect 15640 5056 15646 5073
rect 15663 5056 15669 5073
rect 15640 5039 15669 5056
rect 15640 5022 15646 5039
rect 15663 5022 15669 5039
rect 15640 5005 15669 5022
rect 15640 4988 15646 5005
rect 15663 4988 15669 5005
rect 15640 4980 15669 4988
rect 15684 4980 15705 5080
rect 15720 5073 15749 5080
rect 15720 5056 15726 5073
rect 15743 5056 15749 5073
rect 15720 5039 15749 5056
rect 15720 5022 15726 5039
rect 15743 5022 15749 5039
rect 15720 5005 15749 5022
rect 15720 4988 15726 5005
rect 15743 4988 15749 5005
rect 15720 4980 15749 4988
rect 12450 4433 12479 4440
rect 12450 4416 12456 4433
rect 12473 4416 12479 4433
rect 12450 4399 12479 4416
rect 12450 4382 12456 4399
rect 12473 4382 12479 4399
rect 12450 4365 12479 4382
rect 12450 4348 12456 4365
rect 12473 4348 12479 4365
rect 12450 4340 12479 4348
rect 12494 4340 12515 4440
rect 12530 4433 12559 4440
rect 12530 4416 12536 4433
rect 12553 4416 12559 4433
rect 12530 4399 12559 4416
rect 12530 4382 12536 4399
rect 12553 4382 12559 4399
rect 12530 4365 12559 4382
rect 12530 4348 12536 4365
rect 12553 4348 12559 4365
rect 12530 4340 12559 4348
rect 12574 4433 12603 4440
rect 12574 4416 12580 4433
rect 12597 4416 12603 4433
rect 12574 4399 12603 4416
rect 12574 4382 12580 4399
rect 12597 4382 12603 4399
rect 12574 4365 12603 4382
rect 12574 4348 12580 4365
rect 12597 4348 12603 4365
rect 12574 4340 12603 4348
rect 12618 4433 12647 4440
rect 12618 4416 12624 4433
rect 12641 4416 12647 4433
rect 12618 4399 12647 4416
rect 12618 4382 12624 4399
rect 12641 4382 12647 4399
rect 12618 4365 12647 4382
rect 12618 4348 12624 4365
rect 12641 4348 12647 4365
rect 12618 4340 12647 4348
rect 12662 4340 12683 4440
rect 12698 4433 12727 4440
rect 12698 4416 12704 4433
rect 12721 4416 12727 4433
rect 12698 4399 12727 4416
rect 12698 4382 12704 4399
rect 12721 4382 12727 4399
rect 12698 4365 12727 4382
rect 12698 4348 12704 4365
rect 12721 4348 12727 4365
rect 12698 4340 12727 4348
rect 13061 4433 13090 4440
rect 13061 4416 13067 4433
rect 13084 4416 13090 4433
rect 13061 4399 13090 4416
rect 13061 4382 13067 4399
rect 13084 4382 13090 4399
rect 13061 4365 13090 4382
rect 13061 4348 13067 4365
rect 13084 4348 13090 4365
rect 13061 4340 13090 4348
rect 13105 4340 13126 4440
rect 13141 4433 13170 4440
rect 13141 4416 13147 4433
rect 13164 4416 13170 4433
rect 13141 4399 13170 4416
rect 13141 4382 13147 4399
rect 13164 4382 13170 4399
rect 13141 4365 13170 4382
rect 13141 4348 13147 4365
rect 13164 4348 13170 4365
rect 13141 4340 13170 4348
rect 13185 4433 13214 4440
rect 13185 4416 13191 4433
rect 13208 4416 13214 4433
rect 13185 4399 13214 4416
rect 13185 4382 13191 4399
rect 13208 4382 13214 4399
rect 13185 4365 13214 4382
rect 13185 4348 13191 4365
rect 13208 4348 13214 4365
rect 13185 4340 13214 4348
rect 13229 4433 13258 4440
rect 13229 4416 13235 4433
rect 13252 4416 13258 4433
rect 13229 4399 13258 4416
rect 13229 4382 13235 4399
rect 13252 4382 13258 4399
rect 13229 4365 13258 4382
rect 13229 4348 13235 4365
rect 13252 4348 13258 4365
rect 13229 4340 13258 4348
rect 13273 4340 13294 4440
rect 13309 4433 13338 4440
rect 13309 4416 13315 4433
rect 13332 4416 13338 4433
rect 13309 4399 13338 4416
rect 13309 4382 13315 4399
rect 13332 4382 13338 4399
rect 13309 4365 13338 4382
rect 13309 4348 13315 4365
rect 13332 4348 13338 4365
rect 13309 4340 13338 4348
rect 13672 4433 13701 4440
rect 13672 4416 13678 4433
rect 13695 4416 13701 4433
rect 13672 4399 13701 4416
rect 13672 4382 13678 4399
rect 13695 4382 13701 4399
rect 13672 4365 13701 4382
rect 13672 4348 13678 4365
rect 13695 4348 13701 4365
rect 13672 4340 13701 4348
rect 13716 4340 13737 4440
rect 13752 4433 13781 4440
rect 13752 4416 13758 4433
rect 13775 4416 13781 4433
rect 13752 4399 13781 4416
rect 13752 4382 13758 4399
rect 13775 4382 13781 4399
rect 13752 4365 13781 4382
rect 13752 4348 13758 4365
rect 13775 4348 13781 4365
rect 13752 4340 13781 4348
rect 13796 4433 13825 4440
rect 13796 4416 13802 4433
rect 13819 4416 13825 4433
rect 13796 4399 13825 4416
rect 13796 4382 13802 4399
rect 13819 4382 13825 4399
rect 13796 4365 13825 4382
rect 13796 4348 13802 4365
rect 13819 4348 13825 4365
rect 13796 4340 13825 4348
rect 13840 4433 13869 4440
rect 13840 4416 13846 4433
rect 13863 4416 13869 4433
rect 13840 4399 13869 4416
rect 13840 4382 13846 4399
rect 13863 4382 13869 4399
rect 13840 4365 13869 4382
rect 13840 4348 13846 4365
rect 13863 4348 13869 4365
rect 13840 4340 13869 4348
rect 13884 4340 13905 4440
rect 13920 4433 13949 4440
rect 13920 4416 13926 4433
rect 13943 4416 13949 4433
rect 13920 4399 13949 4416
rect 13920 4382 13926 4399
rect 13943 4382 13949 4399
rect 13920 4365 13949 4382
rect 13920 4348 13926 4365
rect 13943 4348 13949 4365
rect 13920 4340 13949 4348
rect 14250 4433 14279 4440
rect 14250 4416 14256 4433
rect 14273 4416 14279 4433
rect 14250 4399 14279 4416
rect 14250 4382 14256 4399
rect 14273 4382 14279 4399
rect 14250 4365 14279 4382
rect 14250 4348 14256 4365
rect 14273 4348 14279 4365
rect 14250 4340 14279 4348
rect 14294 4340 14315 4440
rect 14330 4433 14359 4440
rect 14330 4416 14336 4433
rect 14353 4416 14359 4433
rect 14330 4399 14359 4416
rect 14330 4382 14336 4399
rect 14353 4382 14359 4399
rect 14330 4365 14359 4382
rect 14330 4348 14336 4365
rect 14353 4348 14359 4365
rect 14330 4340 14359 4348
rect 14374 4433 14403 4440
rect 14374 4416 14380 4433
rect 14397 4416 14403 4433
rect 14374 4399 14403 4416
rect 14374 4382 14380 4399
rect 14397 4382 14403 4399
rect 14374 4365 14403 4382
rect 14374 4348 14380 4365
rect 14397 4348 14403 4365
rect 14374 4340 14403 4348
rect 14418 4433 14447 4440
rect 14418 4416 14424 4433
rect 14441 4416 14447 4433
rect 14418 4399 14447 4416
rect 14418 4382 14424 4399
rect 14441 4382 14447 4399
rect 14418 4365 14447 4382
rect 14418 4348 14424 4365
rect 14441 4348 14447 4365
rect 14418 4340 14447 4348
rect 14462 4340 14483 4440
rect 14498 4433 14527 4440
rect 14498 4416 14504 4433
rect 14521 4416 14527 4433
rect 14498 4399 14527 4416
rect 14498 4382 14504 4399
rect 14521 4382 14527 4399
rect 14498 4365 14527 4382
rect 14498 4348 14504 4365
rect 14521 4348 14527 4365
rect 14498 4340 14527 4348
rect 14861 4433 14890 4440
rect 14861 4416 14867 4433
rect 14884 4416 14890 4433
rect 14861 4399 14890 4416
rect 14861 4382 14867 4399
rect 14884 4382 14890 4399
rect 14861 4365 14890 4382
rect 14861 4348 14867 4365
rect 14884 4348 14890 4365
rect 14861 4340 14890 4348
rect 14905 4340 14926 4440
rect 14941 4433 14970 4440
rect 14941 4416 14947 4433
rect 14964 4416 14970 4433
rect 14941 4399 14970 4416
rect 14941 4382 14947 4399
rect 14964 4382 14970 4399
rect 14941 4365 14970 4382
rect 14941 4348 14947 4365
rect 14964 4348 14970 4365
rect 14941 4340 14970 4348
rect 14985 4433 15014 4440
rect 14985 4416 14991 4433
rect 15008 4416 15014 4433
rect 14985 4399 15014 4416
rect 14985 4382 14991 4399
rect 15008 4382 15014 4399
rect 14985 4365 15014 4382
rect 14985 4348 14991 4365
rect 15008 4348 15014 4365
rect 14985 4340 15014 4348
rect 15029 4433 15058 4440
rect 15029 4416 15035 4433
rect 15052 4416 15058 4433
rect 15029 4399 15058 4416
rect 15029 4382 15035 4399
rect 15052 4382 15058 4399
rect 15029 4365 15058 4382
rect 15029 4348 15035 4365
rect 15052 4348 15058 4365
rect 15029 4340 15058 4348
rect 15073 4340 15094 4440
rect 15109 4433 15138 4440
rect 15109 4416 15115 4433
rect 15132 4416 15138 4433
rect 15109 4399 15138 4416
rect 15109 4382 15115 4399
rect 15132 4382 15138 4399
rect 15109 4365 15138 4382
rect 15109 4348 15115 4365
rect 15132 4348 15138 4365
rect 15109 4340 15138 4348
rect 15472 4433 15501 4440
rect 15472 4416 15478 4433
rect 15495 4416 15501 4433
rect 15472 4399 15501 4416
rect 15472 4382 15478 4399
rect 15495 4382 15501 4399
rect 15472 4365 15501 4382
rect 15472 4348 15478 4365
rect 15495 4348 15501 4365
rect 15472 4340 15501 4348
rect 15516 4340 15537 4440
rect 15552 4433 15581 4440
rect 15552 4416 15558 4433
rect 15575 4416 15581 4433
rect 15552 4399 15581 4416
rect 15552 4382 15558 4399
rect 15575 4382 15581 4399
rect 15552 4365 15581 4382
rect 15552 4348 15558 4365
rect 15575 4348 15581 4365
rect 15552 4340 15581 4348
rect 15596 4433 15625 4440
rect 15596 4416 15602 4433
rect 15619 4416 15625 4433
rect 15596 4399 15625 4416
rect 15596 4382 15602 4399
rect 15619 4382 15625 4399
rect 15596 4365 15625 4382
rect 15596 4348 15602 4365
rect 15619 4348 15625 4365
rect 15596 4340 15625 4348
rect 15640 4433 15669 4440
rect 15640 4416 15646 4433
rect 15663 4416 15669 4433
rect 15640 4399 15669 4416
rect 15640 4382 15646 4399
rect 15663 4382 15669 4399
rect 15640 4365 15669 4382
rect 15640 4348 15646 4365
rect 15663 4348 15669 4365
rect 15640 4340 15669 4348
rect 15684 4340 15705 4440
rect 15720 4433 15749 4440
rect 15720 4416 15726 4433
rect 15743 4416 15749 4433
rect 15720 4399 15749 4416
rect 15720 4382 15726 4399
rect 15743 4382 15749 4399
rect 15720 4365 15749 4382
rect 15720 4348 15726 4365
rect 15743 4348 15749 4365
rect 15720 4340 15749 4348
<< pdiff >>
rect 13141 8039 13170 8044
rect 13141 8022 13147 8039
rect 13164 8022 13170 8039
rect 13141 8005 13170 8022
rect 13141 7988 13147 8005
rect 13164 7988 13170 8005
rect 13141 7971 13170 7988
rect 13141 7954 13147 7971
rect 13164 7954 13170 7971
rect 13141 7937 13170 7954
rect 13141 7920 13147 7937
rect 13164 7920 13170 7937
rect 13141 7903 13170 7920
rect 13141 7886 13147 7903
rect 13164 7886 13170 7903
rect 13141 7869 13170 7886
rect 13141 7852 13147 7869
rect 13164 7852 13170 7869
rect 13141 7844 13170 7852
rect 13185 8039 13214 8044
rect 13185 8022 13191 8039
rect 13208 8022 13214 8039
rect 13185 8005 13214 8022
rect 13185 7988 13191 8005
rect 13208 7988 13214 8005
rect 13185 7971 13214 7988
rect 13185 7954 13191 7971
rect 13208 7954 13214 7971
rect 13185 7937 13214 7954
rect 13185 7920 13191 7937
rect 13208 7920 13214 7937
rect 13185 7903 13214 7920
rect 13185 7886 13191 7903
rect 13208 7886 13214 7903
rect 13185 7869 13214 7886
rect 13185 7852 13191 7869
rect 13208 7852 13214 7869
rect 13185 7844 13214 7852
rect 13229 8039 13258 8044
rect 13229 8022 13235 8039
rect 13252 8022 13258 8039
rect 13229 8005 13258 8022
rect 13229 7988 13235 8005
rect 13252 7988 13258 8005
rect 13229 7971 13258 7988
rect 13229 7954 13235 7971
rect 13252 7954 13258 7971
rect 13229 7937 13258 7954
rect 13229 7920 13235 7937
rect 13252 7920 13258 7937
rect 13229 7903 13258 7920
rect 13229 7886 13235 7903
rect 13252 7886 13258 7903
rect 13229 7869 13258 7886
rect 13229 7852 13235 7869
rect 13252 7852 13258 7869
rect 13229 7844 13258 7852
rect 13752 8039 13781 8044
rect 13752 8022 13758 8039
rect 13775 8022 13781 8039
rect 13752 8005 13781 8022
rect 13752 7988 13758 8005
rect 13775 7988 13781 8005
rect 13752 7971 13781 7988
rect 13752 7954 13758 7971
rect 13775 7954 13781 7971
rect 13752 7937 13781 7954
rect 13752 7920 13758 7937
rect 13775 7920 13781 7937
rect 13752 7903 13781 7920
rect 13752 7886 13758 7903
rect 13775 7886 13781 7903
rect 13752 7869 13781 7886
rect 13752 7852 13758 7869
rect 13775 7852 13781 7869
rect 13752 7844 13781 7852
rect 13796 8039 13825 8044
rect 13796 8022 13802 8039
rect 13819 8022 13825 8039
rect 13796 8005 13825 8022
rect 13796 7988 13802 8005
rect 13819 7988 13825 8005
rect 13796 7971 13825 7988
rect 13796 7954 13802 7971
rect 13819 7954 13825 7971
rect 13796 7937 13825 7954
rect 13796 7920 13802 7937
rect 13819 7920 13825 7937
rect 13796 7903 13825 7920
rect 13796 7886 13802 7903
rect 13819 7886 13825 7903
rect 13796 7869 13825 7886
rect 13796 7852 13802 7869
rect 13819 7852 13825 7869
rect 13796 7844 13825 7852
rect 13840 8039 13869 8044
rect 13840 8022 13846 8039
rect 13863 8022 13869 8039
rect 13840 8005 13869 8022
rect 13840 7988 13846 8005
rect 13863 7988 13869 8005
rect 13840 7971 13869 7988
rect 13840 7954 13846 7971
rect 13863 7954 13869 7971
rect 13840 7937 13869 7954
rect 13840 7920 13846 7937
rect 13863 7920 13869 7937
rect 13840 7903 13869 7920
rect 13840 7886 13846 7903
rect 13863 7886 13869 7903
rect 13840 7869 13869 7886
rect 13840 7852 13846 7869
rect 13863 7852 13869 7869
rect 13840 7844 13869 7852
rect 14330 8039 14359 8044
rect 14330 8022 14336 8039
rect 14353 8022 14359 8039
rect 14330 8005 14359 8022
rect 14330 7988 14336 8005
rect 14353 7988 14359 8005
rect 14330 7971 14359 7988
rect 14330 7954 14336 7971
rect 14353 7954 14359 7971
rect 14330 7937 14359 7954
rect 14330 7920 14336 7937
rect 14353 7920 14359 7937
rect 14330 7903 14359 7920
rect 14330 7886 14336 7903
rect 14353 7886 14359 7903
rect 14330 7869 14359 7886
rect 14330 7852 14336 7869
rect 14353 7852 14359 7869
rect 14330 7844 14359 7852
rect 14374 8039 14403 8044
rect 14374 8022 14380 8039
rect 14397 8022 14403 8039
rect 14374 8005 14403 8022
rect 14374 7988 14380 8005
rect 14397 7988 14403 8005
rect 14374 7971 14403 7988
rect 14374 7954 14380 7971
rect 14397 7954 14403 7971
rect 14374 7937 14403 7954
rect 14374 7920 14380 7937
rect 14397 7920 14403 7937
rect 14374 7903 14403 7920
rect 14374 7886 14380 7903
rect 14397 7886 14403 7903
rect 14374 7869 14403 7886
rect 14374 7852 14380 7869
rect 14397 7852 14403 7869
rect 14374 7844 14403 7852
rect 14418 8039 14447 8044
rect 14418 8022 14424 8039
rect 14441 8022 14447 8039
rect 14418 8005 14447 8022
rect 14418 7988 14424 8005
rect 14441 7988 14447 8005
rect 14418 7971 14447 7988
rect 14418 7954 14424 7971
rect 14441 7954 14447 7971
rect 14418 7937 14447 7954
rect 14418 7920 14424 7937
rect 14441 7920 14447 7937
rect 14418 7903 14447 7920
rect 14418 7886 14424 7903
rect 14441 7886 14447 7903
rect 14418 7869 14447 7886
rect 14418 7852 14424 7869
rect 14441 7852 14447 7869
rect 14418 7844 14447 7852
rect 14941 8039 14970 8044
rect 14941 8022 14947 8039
rect 14964 8022 14970 8039
rect 14941 8005 14970 8022
rect 14941 7988 14947 8005
rect 14964 7988 14970 8005
rect 14941 7971 14970 7988
rect 14941 7954 14947 7971
rect 14964 7954 14970 7971
rect 14941 7937 14970 7954
rect 14941 7920 14947 7937
rect 14964 7920 14970 7937
rect 14941 7903 14970 7920
rect 14941 7886 14947 7903
rect 14964 7886 14970 7903
rect 14941 7869 14970 7886
rect 14941 7852 14947 7869
rect 14964 7852 14970 7869
rect 14941 7844 14970 7852
rect 14985 8039 15014 8044
rect 14985 8022 14991 8039
rect 15008 8022 15014 8039
rect 14985 8005 15014 8022
rect 14985 7988 14991 8005
rect 15008 7988 15014 8005
rect 14985 7971 15014 7988
rect 14985 7954 14991 7971
rect 15008 7954 15014 7971
rect 14985 7937 15014 7954
rect 14985 7920 14991 7937
rect 15008 7920 15014 7937
rect 14985 7903 15014 7920
rect 14985 7886 14991 7903
rect 15008 7886 15014 7903
rect 14985 7869 15014 7886
rect 14985 7852 14991 7869
rect 15008 7852 15014 7869
rect 14985 7844 15014 7852
rect 15029 8039 15058 8044
rect 15029 8022 15035 8039
rect 15052 8022 15058 8039
rect 15029 8005 15058 8022
rect 15029 7988 15035 8005
rect 15052 7988 15058 8005
rect 15029 7971 15058 7988
rect 15029 7954 15035 7971
rect 15052 7954 15058 7971
rect 15029 7937 15058 7954
rect 15029 7920 15035 7937
rect 15052 7920 15058 7937
rect 15029 7903 15058 7920
rect 15029 7886 15035 7903
rect 15052 7886 15058 7903
rect 15029 7869 15058 7886
rect 15029 7852 15035 7869
rect 15052 7852 15058 7869
rect 15029 7844 15058 7852
rect 15552 8039 15581 8044
rect 15552 8022 15558 8039
rect 15575 8022 15581 8039
rect 15552 8005 15581 8022
rect 15552 7988 15558 8005
rect 15575 7988 15581 8005
rect 15552 7971 15581 7988
rect 15552 7954 15558 7971
rect 15575 7954 15581 7971
rect 15552 7937 15581 7954
rect 15552 7920 15558 7937
rect 15575 7920 15581 7937
rect 15552 7903 15581 7920
rect 15552 7886 15558 7903
rect 15575 7886 15581 7903
rect 15552 7869 15581 7886
rect 15552 7852 15558 7869
rect 15575 7852 15581 7869
rect 15552 7844 15581 7852
rect 15596 8039 15625 8044
rect 15596 8022 15602 8039
rect 15619 8022 15625 8039
rect 15596 8005 15625 8022
rect 15596 7988 15602 8005
rect 15619 7988 15625 8005
rect 15596 7971 15625 7988
rect 15596 7954 15602 7971
rect 15619 7954 15625 7971
rect 15596 7937 15625 7954
rect 15596 7920 15602 7937
rect 15619 7920 15625 7937
rect 15596 7903 15625 7920
rect 15596 7886 15602 7903
rect 15619 7886 15625 7903
rect 15596 7869 15625 7886
rect 15596 7852 15602 7869
rect 15619 7852 15625 7869
rect 15596 7844 15625 7852
rect 15640 8039 15669 8044
rect 15640 8022 15646 8039
rect 15663 8022 15669 8039
rect 15640 8005 15669 8022
rect 15640 7988 15646 8005
rect 15663 7988 15669 8005
rect 15640 7971 15669 7988
rect 15640 7954 15646 7971
rect 15663 7954 15669 7971
rect 15640 7937 15669 7954
rect 15640 7920 15646 7937
rect 15663 7920 15669 7937
rect 15640 7903 15669 7920
rect 15640 7886 15646 7903
rect 15663 7886 15669 7903
rect 15640 7869 15669 7886
rect 15640 7852 15646 7869
rect 15663 7852 15669 7869
rect 15640 7844 15669 7852
rect 12530 7389 12559 7394
rect 12530 7372 12536 7389
rect 12553 7372 12559 7389
rect 12530 7355 12559 7372
rect 12530 7338 12536 7355
rect 12553 7338 12559 7355
rect 12530 7321 12559 7338
rect 12530 7304 12536 7321
rect 12553 7304 12559 7321
rect 12530 7287 12559 7304
rect 12530 7270 12536 7287
rect 12553 7270 12559 7287
rect 12530 7253 12559 7270
rect 12530 7236 12536 7253
rect 12553 7236 12559 7253
rect 12530 7219 12559 7236
rect 12530 7202 12536 7219
rect 12553 7202 12559 7219
rect 12530 7194 12559 7202
rect 12574 7389 12603 7394
rect 12574 7372 12580 7389
rect 12597 7372 12603 7389
rect 12574 7355 12603 7372
rect 12574 7338 12580 7355
rect 12597 7338 12603 7355
rect 12574 7321 12603 7338
rect 12574 7304 12580 7321
rect 12597 7304 12603 7321
rect 12574 7287 12603 7304
rect 12574 7270 12580 7287
rect 12597 7270 12603 7287
rect 12574 7253 12603 7270
rect 12574 7236 12580 7253
rect 12597 7236 12603 7253
rect 12574 7219 12603 7236
rect 12574 7202 12580 7219
rect 12597 7202 12603 7219
rect 12574 7194 12603 7202
rect 12618 7389 12647 7394
rect 12618 7372 12624 7389
rect 12641 7372 12647 7389
rect 12618 7355 12647 7372
rect 12618 7338 12624 7355
rect 12641 7338 12647 7355
rect 12618 7321 12647 7338
rect 12618 7304 12624 7321
rect 12641 7304 12647 7321
rect 12618 7287 12647 7304
rect 12618 7270 12624 7287
rect 12641 7270 12647 7287
rect 12618 7253 12647 7270
rect 12618 7236 12624 7253
rect 12641 7236 12647 7253
rect 12618 7219 12647 7236
rect 12618 7202 12624 7219
rect 12641 7202 12647 7219
rect 12618 7194 12647 7202
rect 13141 7389 13170 7394
rect 13141 7372 13147 7389
rect 13164 7372 13170 7389
rect 13141 7355 13170 7372
rect 13141 7338 13147 7355
rect 13164 7338 13170 7355
rect 13141 7321 13170 7338
rect 13141 7304 13147 7321
rect 13164 7304 13170 7321
rect 13141 7287 13170 7304
rect 13141 7270 13147 7287
rect 13164 7270 13170 7287
rect 13141 7253 13170 7270
rect 13141 7236 13147 7253
rect 13164 7236 13170 7253
rect 13141 7219 13170 7236
rect 13141 7202 13147 7219
rect 13164 7202 13170 7219
rect 13141 7194 13170 7202
rect 13185 7389 13214 7394
rect 13185 7372 13191 7389
rect 13208 7372 13214 7389
rect 13185 7355 13214 7372
rect 13185 7338 13191 7355
rect 13208 7338 13214 7355
rect 13185 7321 13214 7338
rect 13185 7304 13191 7321
rect 13208 7304 13214 7321
rect 13185 7287 13214 7304
rect 13185 7270 13191 7287
rect 13208 7270 13214 7287
rect 13185 7253 13214 7270
rect 13185 7236 13191 7253
rect 13208 7236 13214 7253
rect 13185 7219 13214 7236
rect 13185 7202 13191 7219
rect 13208 7202 13214 7219
rect 13185 7194 13214 7202
rect 13229 7389 13258 7394
rect 13229 7372 13235 7389
rect 13252 7372 13258 7389
rect 13229 7355 13258 7372
rect 13229 7338 13235 7355
rect 13252 7338 13258 7355
rect 13229 7321 13258 7338
rect 13229 7304 13235 7321
rect 13252 7304 13258 7321
rect 13229 7287 13258 7304
rect 13229 7270 13235 7287
rect 13252 7270 13258 7287
rect 13229 7253 13258 7270
rect 13229 7236 13235 7253
rect 13252 7236 13258 7253
rect 13229 7219 13258 7236
rect 13229 7202 13235 7219
rect 13252 7202 13258 7219
rect 13229 7194 13258 7202
rect 13752 7389 13781 7394
rect 13752 7372 13758 7389
rect 13775 7372 13781 7389
rect 13752 7355 13781 7372
rect 13752 7338 13758 7355
rect 13775 7338 13781 7355
rect 13752 7321 13781 7338
rect 13752 7304 13758 7321
rect 13775 7304 13781 7321
rect 13752 7287 13781 7304
rect 13752 7270 13758 7287
rect 13775 7270 13781 7287
rect 13752 7253 13781 7270
rect 13752 7236 13758 7253
rect 13775 7236 13781 7253
rect 13752 7219 13781 7236
rect 13752 7202 13758 7219
rect 13775 7202 13781 7219
rect 13752 7194 13781 7202
rect 13796 7389 13825 7394
rect 13796 7372 13802 7389
rect 13819 7372 13825 7389
rect 13796 7355 13825 7372
rect 13796 7338 13802 7355
rect 13819 7338 13825 7355
rect 13796 7321 13825 7338
rect 13796 7304 13802 7321
rect 13819 7304 13825 7321
rect 13796 7287 13825 7304
rect 13796 7270 13802 7287
rect 13819 7270 13825 7287
rect 13796 7253 13825 7270
rect 13796 7236 13802 7253
rect 13819 7236 13825 7253
rect 13796 7219 13825 7236
rect 13796 7202 13802 7219
rect 13819 7202 13825 7219
rect 13796 7194 13825 7202
rect 13840 7389 13869 7394
rect 13840 7372 13846 7389
rect 13863 7372 13869 7389
rect 13840 7355 13869 7372
rect 13840 7338 13846 7355
rect 13863 7338 13869 7355
rect 13840 7321 13869 7338
rect 13840 7304 13846 7321
rect 13863 7304 13869 7321
rect 13840 7287 13869 7304
rect 13840 7270 13846 7287
rect 13863 7270 13869 7287
rect 13840 7253 13869 7270
rect 13840 7236 13846 7253
rect 13863 7236 13869 7253
rect 13840 7219 13869 7236
rect 13840 7202 13846 7219
rect 13863 7202 13869 7219
rect 13840 7194 13869 7202
rect 14330 7389 14359 7394
rect 14330 7372 14336 7389
rect 14353 7372 14359 7389
rect 14330 7355 14359 7372
rect 14330 7338 14336 7355
rect 14353 7338 14359 7355
rect 14330 7321 14359 7338
rect 14330 7304 14336 7321
rect 14353 7304 14359 7321
rect 14330 7287 14359 7304
rect 14330 7270 14336 7287
rect 14353 7270 14359 7287
rect 14330 7253 14359 7270
rect 14330 7236 14336 7253
rect 14353 7236 14359 7253
rect 14330 7219 14359 7236
rect 14330 7202 14336 7219
rect 14353 7202 14359 7219
rect 14330 7194 14359 7202
rect 14374 7389 14403 7394
rect 14374 7372 14380 7389
rect 14397 7372 14403 7389
rect 14374 7355 14403 7372
rect 14374 7338 14380 7355
rect 14397 7338 14403 7355
rect 14374 7321 14403 7338
rect 14374 7304 14380 7321
rect 14397 7304 14403 7321
rect 14374 7287 14403 7304
rect 14374 7270 14380 7287
rect 14397 7270 14403 7287
rect 14374 7253 14403 7270
rect 14374 7236 14380 7253
rect 14397 7236 14403 7253
rect 14374 7219 14403 7236
rect 14374 7202 14380 7219
rect 14397 7202 14403 7219
rect 14374 7194 14403 7202
rect 14418 7389 14447 7394
rect 14418 7372 14424 7389
rect 14441 7372 14447 7389
rect 14418 7355 14447 7372
rect 14418 7338 14424 7355
rect 14441 7338 14447 7355
rect 14418 7321 14447 7338
rect 14418 7304 14424 7321
rect 14441 7304 14447 7321
rect 14418 7287 14447 7304
rect 14418 7270 14424 7287
rect 14441 7270 14447 7287
rect 14418 7253 14447 7270
rect 14418 7236 14424 7253
rect 14441 7236 14447 7253
rect 14418 7219 14447 7236
rect 14418 7202 14424 7219
rect 14441 7202 14447 7219
rect 14418 7194 14447 7202
rect 14941 7389 14970 7394
rect 14941 7372 14947 7389
rect 14964 7372 14970 7389
rect 14941 7355 14970 7372
rect 14941 7338 14947 7355
rect 14964 7338 14970 7355
rect 14941 7321 14970 7338
rect 14941 7304 14947 7321
rect 14964 7304 14970 7321
rect 14941 7287 14970 7304
rect 14941 7270 14947 7287
rect 14964 7270 14970 7287
rect 14941 7253 14970 7270
rect 14941 7236 14947 7253
rect 14964 7236 14970 7253
rect 14941 7219 14970 7236
rect 14941 7202 14947 7219
rect 14964 7202 14970 7219
rect 14941 7194 14970 7202
rect 14985 7389 15014 7394
rect 14985 7372 14991 7389
rect 15008 7372 15014 7389
rect 14985 7355 15014 7372
rect 14985 7338 14991 7355
rect 15008 7338 15014 7355
rect 14985 7321 15014 7338
rect 14985 7304 14991 7321
rect 15008 7304 15014 7321
rect 14985 7287 15014 7304
rect 14985 7270 14991 7287
rect 15008 7270 15014 7287
rect 14985 7253 15014 7270
rect 14985 7236 14991 7253
rect 15008 7236 15014 7253
rect 14985 7219 15014 7236
rect 14985 7202 14991 7219
rect 15008 7202 15014 7219
rect 14985 7194 15014 7202
rect 15029 7389 15058 7394
rect 15029 7372 15035 7389
rect 15052 7372 15058 7389
rect 15029 7355 15058 7372
rect 15029 7338 15035 7355
rect 15052 7338 15058 7355
rect 15029 7321 15058 7338
rect 15029 7304 15035 7321
rect 15052 7304 15058 7321
rect 15029 7287 15058 7304
rect 15029 7270 15035 7287
rect 15052 7270 15058 7287
rect 15029 7253 15058 7270
rect 15029 7236 15035 7253
rect 15052 7236 15058 7253
rect 15029 7219 15058 7236
rect 15029 7202 15035 7219
rect 15052 7202 15058 7219
rect 15029 7194 15058 7202
rect 15552 7389 15581 7394
rect 15552 7372 15558 7389
rect 15575 7372 15581 7389
rect 15552 7355 15581 7372
rect 15552 7338 15558 7355
rect 15575 7338 15581 7355
rect 15552 7321 15581 7338
rect 15552 7304 15558 7321
rect 15575 7304 15581 7321
rect 15552 7287 15581 7304
rect 15552 7270 15558 7287
rect 15575 7270 15581 7287
rect 15552 7253 15581 7270
rect 15552 7236 15558 7253
rect 15575 7236 15581 7253
rect 15552 7219 15581 7236
rect 15552 7202 15558 7219
rect 15575 7202 15581 7219
rect 15552 7194 15581 7202
rect 15596 7389 15625 7394
rect 15596 7372 15602 7389
rect 15619 7372 15625 7389
rect 15596 7355 15625 7372
rect 15596 7338 15602 7355
rect 15619 7338 15625 7355
rect 15596 7321 15625 7338
rect 15596 7304 15602 7321
rect 15619 7304 15625 7321
rect 15596 7287 15625 7304
rect 15596 7270 15602 7287
rect 15619 7270 15625 7287
rect 15596 7253 15625 7270
rect 15596 7236 15602 7253
rect 15619 7236 15625 7253
rect 15596 7219 15625 7236
rect 15596 7202 15602 7219
rect 15619 7202 15625 7219
rect 15596 7194 15625 7202
rect 15640 7389 15669 7394
rect 15640 7372 15646 7389
rect 15663 7372 15669 7389
rect 15640 7355 15669 7372
rect 15640 7338 15646 7355
rect 15663 7338 15669 7355
rect 15640 7321 15669 7338
rect 15640 7304 15646 7321
rect 15663 7304 15669 7321
rect 15640 7287 15669 7304
rect 15640 7270 15646 7287
rect 15663 7270 15669 7287
rect 15640 7253 15669 7270
rect 15640 7236 15646 7253
rect 15663 7236 15669 7253
rect 15640 7219 15669 7236
rect 15640 7202 15646 7219
rect 15663 7202 15669 7219
rect 15640 7194 15669 7202
rect 12530 6749 12559 6754
rect 12530 6732 12536 6749
rect 12553 6732 12559 6749
rect 12530 6715 12559 6732
rect 12530 6698 12536 6715
rect 12553 6698 12559 6715
rect 12530 6681 12559 6698
rect 12530 6664 12536 6681
rect 12553 6664 12559 6681
rect 12530 6647 12559 6664
rect 12530 6630 12536 6647
rect 12553 6630 12559 6647
rect 12530 6613 12559 6630
rect 12530 6596 12536 6613
rect 12553 6596 12559 6613
rect 12530 6579 12559 6596
rect 12530 6562 12536 6579
rect 12553 6562 12559 6579
rect 12530 6554 12559 6562
rect 12574 6749 12603 6754
rect 12574 6732 12580 6749
rect 12597 6732 12603 6749
rect 12574 6715 12603 6732
rect 12574 6698 12580 6715
rect 12597 6698 12603 6715
rect 12574 6681 12603 6698
rect 12574 6664 12580 6681
rect 12597 6664 12603 6681
rect 12574 6647 12603 6664
rect 12574 6630 12580 6647
rect 12597 6630 12603 6647
rect 12574 6613 12603 6630
rect 12574 6596 12580 6613
rect 12597 6596 12603 6613
rect 12574 6579 12603 6596
rect 12574 6562 12580 6579
rect 12597 6562 12603 6579
rect 12574 6554 12603 6562
rect 12618 6749 12647 6754
rect 12618 6732 12624 6749
rect 12641 6732 12647 6749
rect 12618 6715 12647 6732
rect 12618 6698 12624 6715
rect 12641 6698 12647 6715
rect 12618 6681 12647 6698
rect 12618 6664 12624 6681
rect 12641 6664 12647 6681
rect 12618 6647 12647 6664
rect 12618 6630 12624 6647
rect 12641 6630 12647 6647
rect 12618 6613 12647 6630
rect 12618 6596 12624 6613
rect 12641 6596 12647 6613
rect 12618 6579 12647 6596
rect 12618 6562 12624 6579
rect 12641 6562 12647 6579
rect 12618 6554 12647 6562
rect 13141 6749 13170 6754
rect 13141 6732 13147 6749
rect 13164 6732 13170 6749
rect 13141 6715 13170 6732
rect 13141 6698 13147 6715
rect 13164 6698 13170 6715
rect 13141 6681 13170 6698
rect 13141 6664 13147 6681
rect 13164 6664 13170 6681
rect 13141 6647 13170 6664
rect 13141 6630 13147 6647
rect 13164 6630 13170 6647
rect 13141 6613 13170 6630
rect 13141 6596 13147 6613
rect 13164 6596 13170 6613
rect 13141 6579 13170 6596
rect 13141 6562 13147 6579
rect 13164 6562 13170 6579
rect 13141 6554 13170 6562
rect 13185 6749 13214 6754
rect 13185 6732 13191 6749
rect 13208 6732 13214 6749
rect 13185 6715 13214 6732
rect 13185 6698 13191 6715
rect 13208 6698 13214 6715
rect 13185 6681 13214 6698
rect 13185 6664 13191 6681
rect 13208 6664 13214 6681
rect 13185 6647 13214 6664
rect 13185 6630 13191 6647
rect 13208 6630 13214 6647
rect 13185 6613 13214 6630
rect 13185 6596 13191 6613
rect 13208 6596 13214 6613
rect 13185 6579 13214 6596
rect 13185 6562 13191 6579
rect 13208 6562 13214 6579
rect 13185 6554 13214 6562
rect 13229 6749 13258 6754
rect 13229 6732 13235 6749
rect 13252 6732 13258 6749
rect 13229 6715 13258 6732
rect 13229 6698 13235 6715
rect 13252 6698 13258 6715
rect 13229 6681 13258 6698
rect 13229 6664 13235 6681
rect 13252 6664 13258 6681
rect 13229 6647 13258 6664
rect 13229 6630 13235 6647
rect 13252 6630 13258 6647
rect 13229 6613 13258 6630
rect 13229 6596 13235 6613
rect 13252 6596 13258 6613
rect 13229 6579 13258 6596
rect 13229 6562 13235 6579
rect 13252 6562 13258 6579
rect 13229 6554 13258 6562
rect 13752 6749 13781 6754
rect 13752 6732 13758 6749
rect 13775 6732 13781 6749
rect 13752 6715 13781 6732
rect 13752 6698 13758 6715
rect 13775 6698 13781 6715
rect 13752 6681 13781 6698
rect 13752 6664 13758 6681
rect 13775 6664 13781 6681
rect 13752 6647 13781 6664
rect 13752 6630 13758 6647
rect 13775 6630 13781 6647
rect 13752 6613 13781 6630
rect 13752 6596 13758 6613
rect 13775 6596 13781 6613
rect 13752 6579 13781 6596
rect 13752 6562 13758 6579
rect 13775 6562 13781 6579
rect 13752 6554 13781 6562
rect 13796 6749 13825 6754
rect 13796 6732 13802 6749
rect 13819 6732 13825 6749
rect 13796 6715 13825 6732
rect 13796 6698 13802 6715
rect 13819 6698 13825 6715
rect 13796 6681 13825 6698
rect 13796 6664 13802 6681
rect 13819 6664 13825 6681
rect 13796 6647 13825 6664
rect 13796 6630 13802 6647
rect 13819 6630 13825 6647
rect 13796 6613 13825 6630
rect 13796 6596 13802 6613
rect 13819 6596 13825 6613
rect 13796 6579 13825 6596
rect 13796 6562 13802 6579
rect 13819 6562 13825 6579
rect 13796 6554 13825 6562
rect 13840 6749 13869 6754
rect 13840 6732 13846 6749
rect 13863 6732 13869 6749
rect 13840 6715 13869 6732
rect 13840 6698 13846 6715
rect 13863 6698 13869 6715
rect 13840 6681 13869 6698
rect 13840 6664 13846 6681
rect 13863 6664 13869 6681
rect 13840 6647 13869 6664
rect 13840 6630 13846 6647
rect 13863 6630 13869 6647
rect 13840 6613 13869 6630
rect 13840 6596 13846 6613
rect 13863 6596 13869 6613
rect 13840 6579 13869 6596
rect 13840 6562 13846 6579
rect 13863 6562 13869 6579
rect 13840 6554 13869 6562
rect 14330 6749 14359 6754
rect 14330 6732 14336 6749
rect 14353 6732 14359 6749
rect 14330 6715 14359 6732
rect 14330 6698 14336 6715
rect 14353 6698 14359 6715
rect 14330 6681 14359 6698
rect 14330 6664 14336 6681
rect 14353 6664 14359 6681
rect 14330 6647 14359 6664
rect 14330 6630 14336 6647
rect 14353 6630 14359 6647
rect 14330 6613 14359 6630
rect 14330 6596 14336 6613
rect 14353 6596 14359 6613
rect 14330 6579 14359 6596
rect 14330 6562 14336 6579
rect 14353 6562 14359 6579
rect 14330 6554 14359 6562
rect 14374 6749 14403 6754
rect 14374 6732 14380 6749
rect 14397 6732 14403 6749
rect 14374 6715 14403 6732
rect 14374 6698 14380 6715
rect 14397 6698 14403 6715
rect 14374 6681 14403 6698
rect 14374 6664 14380 6681
rect 14397 6664 14403 6681
rect 14374 6647 14403 6664
rect 14374 6630 14380 6647
rect 14397 6630 14403 6647
rect 14374 6613 14403 6630
rect 14374 6596 14380 6613
rect 14397 6596 14403 6613
rect 14374 6579 14403 6596
rect 14374 6562 14380 6579
rect 14397 6562 14403 6579
rect 14374 6554 14403 6562
rect 14418 6749 14447 6754
rect 14418 6732 14424 6749
rect 14441 6732 14447 6749
rect 14418 6715 14447 6732
rect 14418 6698 14424 6715
rect 14441 6698 14447 6715
rect 14418 6681 14447 6698
rect 14418 6664 14424 6681
rect 14441 6664 14447 6681
rect 14418 6647 14447 6664
rect 14418 6630 14424 6647
rect 14441 6630 14447 6647
rect 14418 6613 14447 6630
rect 14418 6596 14424 6613
rect 14441 6596 14447 6613
rect 14418 6579 14447 6596
rect 14418 6562 14424 6579
rect 14441 6562 14447 6579
rect 14418 6554 14447 6562
rect 14941 6749 14970 6754
rect 14941 6732 14947 6749
rect 14964 6732 14970 6749
rect 14941 6715 14970 6732
rect 14941 6698 14947 6715
rect 14964 6698 14970 6715
rect 14941 6681 14970 6698
rect 14941 6664 14947 6681
rect 14964 6664 14970 6681
rect 14941 6647 14970 6664
rect 14941 6630 14947 6647
rect 14964 6630 14970 6647
rect 14941 6613 14970 6630
rect 14941 6596 14947 6613
rect 14964 6596 14970 6613
rect 14941 6579 14970 6596
rect 14941 6562 14947 6579
rect 14964 6562 14970 6579
rect 14941 6554 14970 6562
rect 14985 6749 15014 6754
rect 14985 6732 14991 6749
rect 15008 6732 15014 6749
rect 14985 6715 15014 6732
rect 14985 6698 14991 6715
rect 15008 6698 15014 6715
rect 14985 6681 15014 6698
rect 14985 6664 14991 6681
rect 15008 6664 15014 6681
rect 14985 6647 15014 6664
rect 14985 6630 14991 6647
rect 15008 6630 15014 6647
rect 14985 6613 15014 6630
rect 14985 6596 14991 6613
rect 15008 6596 15014 6613
rect 14985 6579 15014 6596
rect 14985 6562 14991 6579
rect 15008 6562 15014 6579
rect 14985 6554 15014 6562
rect 15029 6749 15058 6754
rect 15029 6732 15035 6749
rect 15052 6732 15058 6749
rect 15029 6715 15058 6732
rect 15029 6698 15035 6715
rect 15052 6698 15058 6715
rect 15029 6681 15058 6698
rect 15029 6664 15035 6681
rect 15052 6664 15058 6681
rect 15029 6647 15058 6664
rect 15029 6630 15035 6647
rect 15052 6630 15058 6647
rect 15029 6613 15058 6630
rect 15029 6596 15035 6613
rect 15052 6596 15058 6613
rect 15029 6579 15058 6596
rect 15029 6562 15035 6579
rect 15052 6562 15058 6579
rect 15029 6554 15058 6562
rect 15552 6749 15581 6754
rect 15552 6732 15558 6749
rect 15575 6732 15581 6749
rect 15552 6715 15581 6732
rect 15552 6698 15558 6715
rect 15575 6698 15581 6715
rect 15552 6681 15581 6698
rect 15552 6664 15558 6681
rect 15575 6664 15581 6681
rect 15552 6647 15581 6664
rect 15552 6630 15558 6647
rect 15575 6630 15581 6647
rect 15552 6613 15581 6630
rect 15552 6596 15558 6613
rect 15575 6596 15581 6613
rect 15552 6579 15581 6596
rect 15552 6562 15558 6579
rect 15575 6562 15581 6579
rect 15552 6554 15581 6562
rect 15596 6749 15625 6754
rect 15596 6732 15602 6749
rect 15619 6732 15625 6749
rect 15596 6715 15625 6732
rect 15596 6698 15602 6715
rect 15619 6698 15625 6715
rect 15596 6681 15625 6698
rect 15596 6664 15602 6681
rect 15619 6664 15625 6681
rect 15596 6647 15625 6664
rect 15596 6630 15602 6647
rect 15619 6630 15625 6647
rect 15596 6613 15625 6630
rect 15596 6596 15602 6613
rect 15619 6596 15625 6613
rect 15596 6579 15625 6596
rect 15596 6562 15602 6579
rect 15619 6562 15625 6579
rect 15596 6554 15625 6562
rect 15640 6749 15669 6754
rect 15640 6732 15646 6749
rect 15663 6732 15669 6749
rect 15640 6715 15669 6732
rect 15640 6698 15646 6715
rect 15663 6698 15669 6715
rect 15640 6681 15669 6698
rect 15640 6664 15646 6681
rect 15663 6664 15669 6681
rect 15640 6647 15669 6664
rect 15640 6630 15646 6647
rect 15663 6630 15669 6647
rect 15640 6613 15669 6630
rect 15640 6596 15646 6613
rect 15663 6596 15669 6613
rect 15640 6579 15669 6596
rect 15640 6562 15646 6579
rect 15663 6562 15669 6579
rect 15640 6554 15669 6562
rect 12530 6099 12559 6104
rect 12530 6082 12536 6099
rect 12553 6082 12559 6099
rect 12530 6065 12559 6082
rect 12530 6048 12536 6065
rect 12553 6048 12559 6065
rect 12530 6031 12559 6048
rect 12530 6014 12536 6031
rect 12553 6014 12559 6031
rect 12530 5997 12559 6014
rect 12530 5980 12536 5997
rect 12553 5980 12559 5997
rect 12530 5963 12559 5980
rect 12530 5946 12536 5963
rect 12553 5946 12559 5963
rect 12530 5929 12559 5946
rect 12530 5912 12536 5929
rect 12553 5912 12559 5929
rect 12530 5904 12559 5912
rect 12574 6099 12603 6104
rect 12574 6082 12580 6099
rect 12597 6082 12603 6099
rect 12574 6065 12603 6082
rect 12574 6048 12580 6065
rect 12597 6048 12603 6065
rect 12574 6031 12603 6048
rect 12574 6014 12580 6031
rect 12597 6014 12603 6031
rect 12574 5997 12603 6014
rect 12574 5980 12580 5997
rect 12597 5980 12603 5997
rect 12574 5963 12603 5980
rect 12574 5946 12580 5963
rect 12597 5946 12603 5963
rect 12574 5929 12603 5946
rect 12574 5912 12580 5929
rect 12597 5912 12603 5929
rect 12574 5904 12603 5912
rect 12618 6099 12647 6104
rect 12618 6082 12624 6099
rect 12641 6082 12647 6099
rect 12618 6065 12647 6082
rect 12618 6048 12624 6065
rect 12641 6048 12647 6065
rect 12618 6031 12647 6048
rect 12618 6014 12624 6031
rect 12641 6014 12647 6031
rect 12618 5997 12647 6014
rect 12618 5980 12624 5997
rect 12641 5980 12647 5997
rect 12618 5963 12647 5980
rect 12618 5946 12624 5963
rect 12641 5946 12647 5963
rect 12618 5929 12647 5946
rect 12618 5912 12624 5929
rect 12641 5912 12647 5929
rect 12618 5904 12647 5912
rect 13141 6099 13170 6104
rect 13141 6082 13147 6099
rect 13164 6082 13170 6099
rect 13141 6065 13170 6082
rect 13141 6048 13147 6065
rect 13164 6048 13170 6065
rect 13141 6031 13170 6048
rect 13141 6014 13147 6031
rect 13164 6014 13170 6031
rect 13141 5997 13170 6014
rect 13141 5980 13147 5997
rect 13164 5980 13170 5997
rect 13141 5963 13170 5980
rect 13141 5946 13147 5963
rect 13164 5946 13170 5963
rect 13141 5929 13170 5946
rect 13141 5912 13147 5929
rect 13164 5912 13170 5929
rect 13141 5904 13170 5912
rect 13185 6099 13214 6104
rect 13185 6082 13191 6099
rect 13208 6082 13214 6099
rect 13185 6065 13214 6082
rect 13185 6048 13191 6065
rect 13208 6048 13214 6065
rect 13185 6031 13214 6048
rect 13185 6014 13191 6031
rect 13208 6014 13214 6031
rect 13185 5997 13214 6014
rect 13185 5980 13191 5997
rect 13208 5980 13214 5997
rect 13185 5963 13214 5980
rect 13185 5946 13191 5963
rect 13208 5946 13214 5963
rect 13185 5929 13214 5946
rect 13185 5912 13191 5929
rect 13208 5912 13214 5929
rect 13185 5904 13214 5912
rect 13229 6099 13258 6104
rect 13229 6082 13235 6099
rect 13252 6082 13258 6099
rect 13229 6065 13258 6082
rect 13229 6048 13235 6065
rect 13252 6048 13258 6065
rect 13229 6031 13258 6048
rect 13229 6014 13235 6031
rect 13252 6014 13258 6031
rect 13229 5997 13258 6014
rect 13229 5980 13235 5997
rect 13252 5980 13258 5997
rect 13229 5963 13258 5980
rect 13229 5946 13235 5963
rect 13252 5946 13258 5963
rect 13229 5929 13258 5946
rect 13229 5912 13235 5929
rect 13252 5912 13258 5929
rect 13229 5904 13258 5912
rect 13752 6099 13781 6104
rect 13752 6082 13758 6099
rect 13775 6082 13781 6099
rect 13752 6065 13781 6082
rect 13752 6048 13758 6065
rect 13775 6048 13781 6065
rect 13752 6031 13781 6048
rect 13752 6014 13758 6031
rect 13775 6014 13781 6031
rect 13752 5997 13781 6014
rect 13752 5980 13758 5997
rect 13775 5980 13781 5997
rect 13752 5963 13781 5980
rect 13752 5946 13758 5963
rect 13775 5946 13781 5963
rect 13752 5929 13781 5946
rect 13752 5912 13758 5929
rect 13775 5912 13781 5929
rect 13752 5904 13781 5912
rect 13796 6099 13825 6104
rect 13796 6082 13802 6099
rect 13819 6082 13825 6099
rect 13796 6065 13825 6082
rect 13796 6048 13802 6065
rect 13819 6048 13825 6065
rect 13796 6031 13825 6048
rect 13796 6014 13802 6031
rect 13819 6014 13825 6031
rect 13796 5997 13825 6014
rect 13796 5980 13802 5997
rect 13819 5980 13825 5997
rect 13796 5963 13825 5980
rect 13796 5946 13802 5963
rect 13819 5946 13825 5963
rect 13796 5929 13825 5946
rect 13796 5912 13802 5929
rect 13819 5912 13825 5929
rect 13796 5904 13825 5912
rect 13840 6099 13869 6104
rect 13840 6082 13846 6099
rect 13863 6082 13869 6099
rect 13840 6065 13869 6082
rect 13840 6048 13846 6065
rect 13863 6048 13869 6065
rect 13840 6031 13869 6048
rect 13840 6014 13846 6031
rect 13863 6014 13869 6031
rect 13840 5997 13869 6014
rect 13840 5980 13846 5997
rect 13863 5980 13869 5997
rect 13840 5963 13869 5980
rect 13840 5946 13846 5963
rect 13863 5946 13869 5963
rect 13840 5929 13869 5946
rect 13840 5912 13846 5929
rect 13863 5912 13869 5929
rect 13840 5904 13869 5912
rect 14330 6099 14359 6104
rect 14330 6082 14336 6099
rect 14353 6082 14359 6099
rect 14330 6065 14359 6082
rect 14330 6048 14336 6065
rect 14353 6048 14359 6065
rect 14330 6031 14359 6048
rect 14330 6014 14336 6031
rect 14353 6014 14359 6031
rect 14330 5997 14359 6014
rect 14330 5980 14336 5997
rect 14353 5980 14359 5997
rect 14330 5963 14359 5980
rect 14330 5946 14336 5963
rect 14353 5946 14359 5963
rect 14330 5929 14359 5946
rect 14330 5912 14336 5929
rect 14353 5912 14359 5929
rect 14330 5904 14359 5912
rect 14374 6099 14403 6104
rect 14374 6082 14380 6099
rect 14397 6082 14403 6099
rect 14374 6065 14403 6082
rect 14374 6048 14380 6065
rect 14397 6048 14403 6065
rect 14374 6031 14403 6048
rect 14374 6014 14380 6031
rect 14397 6014 14403 6031
rect 14374 5997 14403 6014
rect 14374 5980 14380 5997
rect 14397 5980 14403 5997
rect 14374 5963 14403 5980
rect 14374 5946 14380 5963
rect 14397 5946 14403 5963
rect 14374 5929 14403 5946
rect 14374 5912 14380 5929
rect 14397 5912 14403 5929
rect 14374 5904 14403 5912
rect 14418 6099 14447 6104
rect 14418 6082 14424 6099
rect 14441 6082 14447 6099
rect 14418 6065 14447 6082
rect 14418 6048 14424 6065
rect 14441 6048 14447 6065
rect 14418 6031 14447 6048
rect 14418 6014 14424 6031
rect 14441 6014 14447 6031
rect 14418 5997 14447 6014
rect 14418 5980 14424 5997
rect 14441 5980 14447 5997
rect 14418 5963 14447 5980
rect 14418 5946 14424 5963
rect 14441 5946 14447 5963
rect 14418 5929 14447 5946
rect 14418 5912 14424 5929
rect 14441 5912 14447 5929
rect 14418 5904 14447 5912
rect 14941 6099 14970 6104
rect 14941 6082 14947 6099
rect 14964 6082 14970 6099
rect 14941 6065 14970 6082
rect 14941 6048 14947 6065
rect 14964 6048 14970 6065
rect 14941 6031 14970 6048
rect 14941 6014 14947 6031
rect 14964 6014 14970 6031
rect 14941 5997 14970 6014
rect 14941 5980 14947 5997
rect 14964 5980 14970 5997
rect 14941 5963 14970 5980
rect 14941 5946 14947 5963
rect 14964 5946 14970 5963
rect 14941 5929 14970 5946
rect 14941 5912 14947 5929
rect 14964 5912 14970 5929
rect 14941 5904 14970 5912
rect 14985 6099 15014 6104
rect 14985 6082 14991 6099
rect 15008 6082 15014 6099
rect 14985 6065 15014 6082
rect 14985 6048 14991 6065
rect 15008 6048 15014 6065
rect 14985 6031 15014 6048
rect 14985 6014 14991 6031
rect 15008 6014 15014 6031
rect 14985 5997 15014 6014
rect 14985 5980 14991 5997
rect 15008 5980 15014 5997
rect 14985 5963 15014 5980
rect 14985 5946 14991 5963
rect 15008 5946 15014 5963
rect 14985 5929 15014 5946
rect 14985 5912 14991 5929
rect 15008 5912 15014 5929
rect 14985 5904 15014 5912
rect 15029 6099 15058 6104
rect 15029 6082 15035 6099
rect 15052 6082 15058 6099
rect 15029 6065 15058 6082
rect 15029 6048 15035 6065
rect 15052 6048 15058 6065
rect 15029 6031 15058 6048
rect 15029 6014 15035 6031
rect 15052 6014 15058 6031
rect 15029 5997 15058 6014
rect 15029 5980 15035 5997
rect 15052 5980 15058 5997
rect 15029 5963 15058 5980
rect 15029 5946 15035 5963
rect 15052 5946 15058 5963
rect 15029 5929 15058 5946
rect 15029 5912 15035 5929
rect 15052 5912 15058 5929
rect 15029 5904 15058 5912
rect 15552 6099 15581 6104
rect 15552 6082 15558 6099
rect 15575 6082 15581 6099
rect 15552 6065 15581 6082
rect 15552 6048 15558 6065
rect 15575 6048 15581 6065
rect 15552 6031 15581 6048
rect 15552 6014 15558 6031
rect 15575 6014 15581 6031
rect 15552 5997 15581 6014
rect 15552 5980 15558 5997
rect 15575 5980 15581 5997
rect 15552 5963 15581 5980
rect 15552 5946 15558 5963
rect 15575 5946 15581 5963
rect 15552 5929 15581 5946
rect 15552 5912 15558 5929
rect 15575 5912 15581 5929
rect 15552 5904 15581 5912
rect 15596 6099 15625 6104
rect 15596 6082 15602 6099
rect 15619 6082 15625 6099
rect 15596 6065 15625 6082
rect 15596 6048 15602 6065
rect 15619 6048 15625 6065
rect 15596 6031 15625 6048
rect 15596 6014 15602 6031
rect 15619 6014 15625 6031
rect 15596 5997 15625 6014
rect 15596 5980 15602 5997
rect 15619 5980 15625 5997
rect 15596 5963 15625 5980
rect 15596 5946 15602 5963
rect 15619 5946 15625 5963
rect 15596 5929 15625 5946
rect 15596 5912 15602 5929
rect 15619 5912 15625 5929
rect 15596 5904 15625 5912
rect 15640 6099 15669 6104
rect 15640 6082 15646 6099
rect 15663 6082 15669 6099
rect 15640 6065 15669 6082
rect 15640 6048 15646 6065
rect 15663 6048 15669 6065
rect 15640 6031 15669 6048
rect 15640 6014 15646 6031
rect 15663 6014 15669 6031
rect 15640 5997 15669 6014
rect 15640 5980 15646 5997
rect 15663 5980 15669 5997
rect 15640 5963 15669 5980
rect 15640 5946 15646 5963
rect 15663 5946 15669 5963
rect 15640 5929 15669 5946
rect 15640 5912 15646 5929
rect 15663 5912 15669 5929
rect 15640 5904 15669 5912
rect 12530 5449 12559 5454
rect 12530 5432 12536 5449
rect 12553 5432 12559 5449
rect 12530 5415 12559 5432
rect 12530 5398 12536 5415
rect 12553 5398 12559 5415
rect 12530 5381 12559 5398
rect 12530 5364 12536 5381
rect 12553 5364 12559 5381
rect 12530 5347 12559 5364
rect 12530 5330 12536 5347
rect 12553 5330 12559 5347
rect 12530 5313 12559 5330
rect 12530 5296 12536 5313
rect 12553 5296 12559 5313
rect 12530 5279 12559 5296
rect 12530 5262 12536 5279
rect 12553 5262 12559 5279
rect 12530 5254 12559 5262
rect 12574 5449 12603 5454
rect 12574 5432 12580 5449
rect 12597 5432 12603 5449
rect 12574 5415 12603 5432
rect 12574 5398 12580 5415
rect 12597 5398 12603 5415
rect 12574 5381 12603 5398
rect 12574 5364 12580 5381
rect 12597 5364 12603 5381
rect 12574 5347 12603 5364
rect 12574 5330 12580 5347
rect 12597 5330 12603 5347
rect 12574 5313 12603 5330
rect 12574 5296 12580 5313
rect 12597 5296 12603 5313
rect 12574 5279 12603 5296
rect 12574 5262 12580 5279
rect 12597 5262 12603 5279
rect 12574 5254 12603 5262
rect 12618 5449 12647 5454
rect 12618 5432 12624 5449
rect 12641 5432 12647 5449
rect 12618 5415 12647 5432
rect 12618 5398 12624 5415
rect 12641 5398 12647 5415
rect 12618 5381 12647 5398
rect 12618 5364 12624 5381
rect 12641 5364 12647 5381
rect 12618 5347 12647 5364
rect 12618 5330 12624 5347
rect 12641 5330 12647 5347
rect 12618 5313 12647 5330
rect 12618 5296 12624 5313
rect 12641 5296 12647 5313
rect 12618 5279 12647 5296
rect 12618 5262 12624 5279
rect 12641 5262 12647 5279
rect 12618 5254 12647 5262
rect 13141 5449 13170 5454
rect 13141 5432 13147 5449
rect 13164 5432 13170 5449
rect 13141 5415 13170 5432
rect 13141 5398 13147 5415
rect 13164 5398 13170 5415
rect 13141 5381 13170 5398
rect 13141 5364 13147 5381
rect 13164 5364 13170 5381
rect 13141 5347 13170 5364
rect 13141 5330 13147 5347
rect 13164 5330 13170 5347
rect 13141 5313 13170 5330
rect 13141 5296 13147 5313
rect 13164 5296 13170 5313
rect 13141 5279 13170 5296
rect 13141 5262 13147 5279
rect 13164 5262 13170 5279
rect 13141 5254 13170 5262
rect 13185 5449 13214 5454
rect 13185 5432 13191 5449
rect 13208 5432 13214 5449
rect 13185 5415 13214 5432
rect 13185 5398 13191 5415
rect 13208 5398 13214 5415
rect 13185 5381 13214 5398
rect 13185 5364 13191 5381
rect 13208 5364 13214 5381
rect 13185 5347 13214 5364
rect 13185 5330 13191 5347
rect 13208 5330 13214 5347
rect 13185 5313 13214 5330
rect 13185 5296 13191 5313
rect 13208 5296 13214 5313
rect 13185 5279 13214 5296
rect 13185 5262 13191 5279
rect 13208 5262 13214 5279
rect 13185 5254 13214 5262
rect 13229 5449 13258 5454
rect 13229 5432 13235 5449
rect 13252 5432 13258 5449
rect 13229 5415 13258 5432
rect 13229 5398 13235 5415
rect 13252 5398 13258 5415
rect 13229 5381 13258 5398
rect 13229 5364 13235 5381
rect 13252 5364 13258 5381
rect 13229 5347 13258 5364
rect 13229 5330 13235 5347
rect 13252 5330 13258 5347
rect 13229 5313 13258 5330
rect 13229 5296 13235 5313
rect 13252 5296 13258 5313
rect 13229 5279 13258 5296
rect 13229 5262 13235 5279
rect 13252 5262 13258 5279
rect 13229 5254 13258 5262
rect 13752 5449 13781 5454
rect 13752 5432 13758 5449
rect 13775 5432 13781 5449
rect 13752 5415 13781 5432
rect 13752 5398 13758 5415
rect 13775 5398 13781 5415
rect 13752 5381 13781 5398
rect 13752 5364 13758 5381
rect 13775 5364 13781 5381
rect 13752 5347 13781 5364
rect 13752 5330 13758 5347
rect 13775 5330 13781 5347
rect 13752 5313 13781 5330
rect 13752 5296 13758 5313
rect 13775 5296 13781 5313
rect 13752 5279 13781 5296
rect 13752 5262 13758 5279
rect 13775 5262 13781 5279
rect 13752 5254 13781 5262
rect 13796 5449 13825 5454
rect 13796 5432 13802 5449
rect 13819 5432 13825 5449
rect 13796 5415 13825 5432
rect 13796 5398 13802 5415
rect 13819 5398 13825 5415
rect 13796 5381 13825 5398
rect 13796 5364 13802 5381
rect 13819 5364 13825 5381
rect 13796 5347 13825 5364
rect 13796 5330 13802 5347
rect 13819 5330 13825 5347
rect 13796 5313 13825 5330
rect 13796 5296 13802 5313
rect 13819 5296 13825 5313
rect 13796 5279 13825 5296
rect 13796 5262 13802 5279
rect 13819 5262 13825 5279
rect 13796 5254 13825 5262
rect 13840 5449 13869 5454
rect 13840 5432 13846 5449
rect 13863 5432 13869 5449
rect 13840 5415 13869 5432
rect 13840 5398 13846 5415
rect 13863 5398 13869 5415
rect 13840 5381 13869 5398
rect 13840 5364 13846 5381
rect 13863 5364 13869 5381
rect 13840 5347 13869 5364
rect 13840 5330 13846 5347
rect 13863 5330 13869 5347
rect 13840 5313 13869 5330
rect 13840 5296 13846 5313
rect 13863 5296 13869 5313
rect 13840 5279 13869 5296
rect 13840 5262 13846 5279
rect 13863 5262 13869 5279
rect 13840 5254 13869 5262
rect 14330 5449 14359 5454
rect 14330 5432 14336 5449
rect 14353 5432 14359 5449
rect 14330 5415 14359 5432
rect 14330 5398 14336 5415
rect 14353 5398 14359 5415
rect 14330 5381 14359 5398
rect 14330 5364 14336 5381
rect 14353 5364 14359 5381
rect 14330 5347 14359 5364
rect 14330 5330 14336 5347
rect 14353 5330 14359 5347
rect 14330 5313 14359 5330
rect 14330 5296 14336 5313
rect 14353 5296 14359 5313
rect 14330 5279 14359 5296
rect 14330 5262 14336 5279
rect 14353 5262 14359 5279
rect 14330 5254 14359 5262
rect 14374 5449 14403 5454
rect 14374 5432 14380 5449
rect 14397 5432 14403 5449
rect 14374 5415 14403 5432
rect 14374 5398 14380 5415
rect 14397 5398 14403 5415
rect 14374 5381 14403 5398
rect 14374 5364 14380 5381
rect 14397 5364 14403 5381
rect 14374 5347 14403 5364
rect 14374 5330 14380 5347
rect 14397 5330 14403 5347
rect 14374 5313 14403 5330
rect 14374 5296 14380 5313
rect 14397 5296 14403 5313
rect 14374 5279 14403 5296
rect 14374 5262 14380 5279
rect 14397 5262 14403 5279
rect 14374 5254 14403 5262
rect 14418 5449 14447 5454
rect 14418 5432 14424 5449
rect 14441 5432 14447 5449
rect 14418 5415 14447 5432
rect 14418 5398 14424 5415
rect 14441 5398 14447 5415
rect 14418 5381 14447 5398
rect 14418 5364 14424 5381
rect 14441 5364 14447 5381
rect 14418 5347 14447 5364
rect 14418 5330 14424 5347
rect 14441 5330 14447 5347
rect 14418 5313 14447 5330
rect 14418 5296 14424 5313
rect 14441 5296 14447 5313
rect 14418 5279 14447 5296
rect 14418 5262 14424 5279
rect 14441 5262 14447 5279
rect 14418 5254 14447 5262
rect 14941 5449 14970 5454
rect 14941 5432 14947 5449
rect 14964 5432 14970 5449
rect 14941 5415 14970 5432
rect 14941 5398 14947 5415
rect 14964 5398 14970 5415
rect 14941 5381 14970 5398
rect 14941 5364 14947 5381
rect 14964 5364 14970 5381
rect 14941 5347 14970 5364
rect 14941 5330 14947 5347
rect 14964 5330 14970 5347
rect 14941 5313 14970 5330
rect 14941 5296 14947 5313
rect 14964 5296 14970 5313
rect 14941 5279 14970 5296
rect 14941 5262 14947 5279
rect 14964 5262 14970 5279
rect 14941 5254 14970 5262
rect 14985 5449 15014 5454
rect 14985 5432 14991 5449
rect 15008 5432 15014 5449
rect 14985 5415 15014 5432
rect 14985 5398 14991 5415
rect 15008 5398 15014 5415
rect 14985 5381 15014 5398
rect 14985 5364 14991 5381
rect 15008 5364 15014 5381
rect 14985 5347 15014 5364
rect 14985 5330 14991 5347
rect 15008 5330 15014 5347
rect 14985 5313 15014 5330
rect 14985 5296 14991 5313
rect 15008 5296 15014 5313
rect 14985 5279 15014 5296
rect 14985 5262 14991 5279
rect 15008 5262 15014 5279
rect 14985 5254 15014 5262
rect 15029 5449 15058 5454
rect 15029 5432 15035 5449
rect 15052 5432 15058 5449
rect 15029 5415 15058 5432
rect 15029 5398 15035 5415
rect 15052 5398 15058 5415
rect 15029 5381 15058 5398
rect 15029 5364 15035 5381
rect 15052 5364 15058 5381
rect 15029 5347 15058 5364
rect 15029 5330 15035 5347
rect 15052 5330 15058 5347
rect 15029 5313 15058 5330
rect 15029 5296 15035 5313
rect 15052 5296 15058 5313
rect 15029 5279 15058 5296
rect 15029 5262 15035 5279
rect 15052 5262 15058 5279
rect 15029 5254 15058 5262
rect 15552 5449 15581 5454
rect 15552 5432 15558 5449
rect 15575 5432 15581 5449
rect 15552 5415 15581 5432
rect 15552 5398 15558 5415
rect 15575 5398 15581 5415
rect 15552 5381 15581 5398
rect 15552 5364 15558 5381
rect 15575 5364 15581 5381
rect 15552 5347 15581 5364
rect 15552 5330 15558 5347
rect 15575 5330 15581 5347
rect 15552 5313 15581 5330
rect 15552 5296 15558 5313
rect 15575 5296 15581 5313
rect 15552 5279 15581 5296
rect 15552 5262 15558 5279
rect 15575 5262 15581 5279
rect 15552 5254 15581 5262
rect 15596 5449 15625 5454
rect 15596 5432 15602 5449
rect 15619 5432 15625 5449
rect 15596 5415 15625 5432
rect 15596 5398 15602 5415
rect 15619 5398 15625 5415
rect 15596 5381 15625 5398
rect 15596 5364 15602 5381
rect 15619 5364 15625 5381
rect 15596 5347 15625 5364
rect 15596 5330 15602 5347
rect 15619 5330 15625 5347
rect 15596 5313 15625 5330
rect 15596 5296 15602 5313
rect 15619 5296 15625 5313
rect 15596 5279 15625 5296
rect 15596 5262 15602 5279
rect 15619 5262 15625 5279
rect 15596 5254 15625 5262
rect 15640 5449 15669 5454
rect 15640 5432 15646 5449
rect 15663 5432 15669 5449
rect 15640 5415 15669 5432
rect 15640 5398 15646 5415
rect 15663 5398 15669 5415
rect 15640 5381 15669 5398
rect 15640 5364 15646 5381
rect 15663 5364 15669 5381
rect 15640 5347 15669 5364
rect 15640 5330 15646 5347
rect 15663 5330 15669 5347
rect 15640 5313 15669 5330
rect 15640 5296 15646 5313
rect 15663 5296 15669 5313
rect 15640 5279 15669 5296
rect 15640 5262 15646 5279
rect 15663 5262 15669 5279
rect 15640 5254 15669 5262
rect 12530 4809 12559 4814
rect 12530 4792 12536 4809
rect 12553 4792 12559 4809
rect 12530 4775 12559 4792
rect 12530 4758 12536 4775
rect 12553 4758 12559 4775
rect 12530 4741 12559 4758
rect 12530 4724 12536 4741
rect 12553 4724 12559 4741
rect 12530 4707 12559 4724
rect 12530 4690 12536 4707
rect 12553 4690 12559 4707
rect 12530 4673 12559 4690
rect 12530 4656 12536 4673
rect 12553 4656 12559 4673
rect 12530 4639 12559 4656
rect 12530 4622 12536 4639
rect 12553 4622 12559 4639
rect 12530 4614 12559 4622
rect 12574 4809 12603 4814
rect 12574 4792 12580 4809
rect 12597 4792 12603 4809
rect 12574 4775 12603 4792
rect 12574 4758 12580 4775
rect 12597 4758 12603 4775
rect 12574 4741 12603 4758
rect 12574 4724 12580 4741
rect 12597 4724 12603 4741
rect 12574 4707 12603 4724
rect 12574 4690 12580 4707
rect 12597 4690 12603 4707
rect 12574 4673 12603 4690
rect 12574 4656 12580 4673
rect 12597 4656 12603 4673
rect 12574 4639 12603 4656
rect 12574 4622 12580 4639
rect 12597 4622 12603 4639
rect 12574 4614 12603 4622
rect 12618 4809 12647 4814
rect 12618 4792 12624 4809
rect 12641 4792 12647 4809
rect 12618 4775 12647 4792
rect 12618 4758 12624 4775
rect 12641 4758 12647 4775
rect 12618 4741 12647 4758
rect 12618 4724 12624 4741
rect 12641 4724 12647 4741
rect 12618 4707 12647 4724
rect 12618 4690 12624 4707
rect 12641 4690 12647 4707
rect 12618 4673 12647 4690
rect 12618 4656 12624 4673
rect 12641 4656 12647 4673
rect 12618 4639 12647 4656
rect 12618 4622 12624 4639
rect 12641 4622 12647 4639
rect 12618 4614 12647 4622
rect 13141 4809 13170 4814
rect 13141 4792 13147 4809
rect 13164 4792 13170 4809
rect 13141 4775 13170 4792
rect 13141 4758 13147 4775
rect 13164 4758 13170 4775
rect 13141 4741 13170 4758
rect 13141 4724 13147 4741
rect 13164 4724 13170 4741
rect 13141 4707 13170 4724
rect 13141 4690 13147 4707
rect 13164 4690 13170 4707
rect 13141 4673 13170 4690
rect 13141 4656 13147 4673
rect 13164 4656 13170 4673
rect 13141 4639 13170 4656
rect 13141 4622 13147 4639
rect 13164 4622 13170 4639
rect 13141 4614 13170 4622
rect 13185 4809 13214 4814
rect 13185 4792 13191 4809
rect 13208 4792 13214 4809
rect 13185 4775 13214 4792
rect 13185 4758 13191 4775
rect 13208 4758 13214 4775
rect 13185 4741 13214 4758
rect 13185 4724 13191 4741
rect 13208 4724 13214 4741
rect 13185 4707 13214 4724
rect 13185 4690 13191 4707
rect 13208 4690 13214 4707
rect 13185 4673 13214 4690
rect 13185 4656 13191 4673
rect 13208 4656 13214 4673
rect 13185 4639 13214 4656
rect 13185 4622 13191 4639
rect 13208 4622 13214 4639
rect 13185 4614 13214 4622
rect 13229 4809 13258 4814
rect 13229 4792 13235 4809
rect 13252 4792 13258 4809
rect 13229 4775 13258 4792
rect 13229 4758 13235 4775
rect 13252 4758 13258 4775
rect 13229 4741 13258 4758
rect 13229 4724 13235 4741
rect 13252 4724 13258 4741
rect 13229 4707 13258 4724
rect 13229 4690 13235 4707
rect 13252 4690 13258 4707
rect 13229 4673 13258 4690
rect 13229 4656 13235 4673
rect 13252 4656 13258 4673
rect 13229 4639 13258 4656
rect 13229 4622 13235 4639
rect 13252 4622 13258 4639
rect 13229 4614 13258 4622
rect 13752 4809 13781 4814
rect 13752 4792 13758 4809
rect 13775 4792 13781 4809
rect 13752 4775 13781 4792
rect 13752 4758 13758 4775
rect 13775 4758 13781 4775
rect 13752 4741 13781 4758
rect 13752 4724 13758 4741
rect 13775 4724 13781 4741
rect 13752 4707 13781 4724
rect 13752 4690 13758 4707
rect 13775 4690 13781 4707
rect 13752 4673 13781 4690
rect 13752 4656 13758 4673
rect 13775 4656 13781 4673
rect 13752 4639 13781 4656
rect 13752 4622 13758 4639
rect 13775 4622 13781 4639
rect 13752 4614 13781 4622
rect 13796 4809 13825 4814
rect 13796 4792 13802 4809
rect 13819 4792 13825 4809
rect 13796 4775 13825 4792
rect 13796 4758 13802 4775
rect 13819 4758 13825 4775
rect 13796 4741 13825 4758
rect 13796 4724 13802 4741
rect 13819 4724 13825 4741
rect 13796 4707 13825 4724
rect 13796 4690 13802 4707
rect 13819 4690 13825 4707
rect 13796 4673 13825 4690
rect 13796 4656 13802 4673
rect 13819 4656 13825 4673
rect 13796 4639 13825 4656
rect 13796 4622 13802 4639
rect 13819 4622 13825 4639
rect 13796 4614 13825 4622
rect 13840 4809 13869 4814
rect 13840 4792 13846 4809
rect 13863 4792 13869 4809
rect 13840 4775 13869 4792
rect 13840 4758 13846 4775
rect 13863 4758 13869 4775
rect 13840 4741 13869 4758
rect 13840 4724 13846 4741
rect 13863 4724 13869 4741
rect 13840 4707 13869 4724
rect 13840 4690 13846 4707
rect 13863 4690 13869 4707
rect 13840 4673 13869 4690
rect 13840 4656 13846 4673
rect 13863 4656 13869 4673
rect 13840 4639 13869 4656
rect 13840 4622 13846 4639
rect 13863 4622 13869 4639
rect 13840 4614 13869 4622
rect 14330 4809 14359 4814
rect 14330 4792 14336 4809
rect 14353 4792 14359 4809
rect 14330 4775 14359 4792
rect 14330 4758 14336 4775
rect 14353 4758 14359 4775
rect 14330 4741 14359 4758
rect 14330 4724 14336 4741
rect 14353 4724 14359 4741
rect 14330 4707 14359 4724
rect 14330 4690 14336 4707
rect 14353 4690 14359 4707
rect 14330 4673 14359 4690
rect 14330 4656 14336 4673
rect 14353 4656 14359 4673
rect 14330 4639 14359 4656
rect 14330 4622 14336 4639
rect 14353 4622 14359 4639
rect 14330 4614 14359 4622
rect 14374 4809 14403 4814
rect 14374 4792 14380 4809
rect 14397 4792 14403 4809
rect 14374 4775 14403 4792
rect 14374 4758 14380 4775
rect 14397 4758 14403 4775
rect 14374 4741 14403 4758
rect 14374 4724 14380 4741
rect 14397 4724 14403 4741
rect 14374 4707 14403 4724
rect 14374 4690 14380 4707
rect 14397 4690 14403 4707
rect 14374 4673 14403 4690
rect 14374 4656 14380 4673
rect 14397 4656 14403 4673
rect 14374 4639 14403 4656
rect 14374 4622 14380 4639
rect 14397 4622 14403 4639
rect 14374 4614 14403 4622
rect 14418 4809 14447 4814
rect 14418 4792 14424 4809
rect 14441 4792 14447 4809
rect 14418 4775 14447 4792
rect 14418 4758 14424 4775
rect 14441 4758 14447 4775
rect 14418 4741 14447 4758
rect 14418 4724 14424 4741
rect 14441 4724 14447 4741
rect 14418 4707 14447 4724
rect 14418 4690 14424 4707
rect 14441 4690 14447 4707
rect 14418 4673 14447 4690
rect 14418 4656 14424 4673
rect 14441 4656 14447 4673
rect 14418 4639 14447 4656
rect 14418 4622 14424 4639
rect 14441 4622 14447 4639
rect 14418 4614 14447 4622
rect 14941 4809 14970 4814
rect 14941 4792 14947 4809
rect 14964 4792 14970 4809
rect 14941 4775 14970 4792
rect 14941 4758 14947 4775
rect 14964 4758 14970 4775
rect 14941 4741 14970 4758
rect 14941 4724 14947 4741
rect 14964 4724 14970 4741
rect 14941 4707 14970 4724
rect 14941 4690 14947 4707
rect 14964 4690 14970 4707
rect 14941 4673 14970 4690
rect 14941 4656 14947 4673
rect 14964 4656 14970 4673
rect 14941 4639 14970 4656
rect 14941 4622 14947 4639
rect 14964 4622 14970 4639
rect 14941 4614 14970 4622
rect 14985 4809 15014 4814
rect 14985 4792 14991 4809
rect 15008 4792 15014 4809
rect 14985 4775 15014 4792
rect 14985 4758 14991 4775
rect 15008 4758 15014 4775
rect 14985 4741 15014 4758
rect 14985 4724 14991 4741
rect 15008 4724 15014 4741
rect 14985 4707 15014 4724
rect 14985 4690 14991 4707
rect 15008 4690 15014 4707
rect 14985 4673 15014 4690
rect 14985 4656 14991 4673
rect 15008 4656 15014 4673
rect 14985 4639 15014 4656
rect 14985 4622 14991 4639
rect 15008 4622 15014 4639
rect 14985 4614 15014 4622
rect 15029 4809 15058 4814
rect 15029 4792 15035 4809
rect 15052 4792 15058 4809
rect 15029 4775 15058 4792
rect 15029 4758 15035 4775
rect 15052 4758 15058 4775
rect 15029 4741 15058 4758
rect 15029 4724 15035 4741
rect 15052 4724 15058 4741
rect 15029 4707 15058 4724
rect 15029 4690 15035 4707
rect 15052 4690 15058 4707
rect 15029 4673 15058 4690
rect 15029 4656 15035 4673
rect 15052 4656 15058 4673
rect 15029 4639 15058 4656
rect 15029 4622 15035 4639
rect 15052 4622 15058 4639
rect 15029 4614 15058 4622
rect 15552 4809 15581 4814
rect 15552 4792 15558 4809
rect 15575 4792 15581 4809
rect 15552 4775 15581 4792
rect 15552 4758 15558 4775
rect 15575 4758 15581 4775
rect 15552 4741 15581 4758
rect 15552 4724 15558 4741
rect 15575 4724 15581 4741
rect 15552 4707 15581 4724
rect 15552 4690 15558 4707
rect 15575 4690 15581 4707
rect 15552 4673 15581 4690
rect 15552 4656 15558 4673
rect 15575 4656 15581 4673
rect 15552 4639 15581 4656
rect 15552 4622 15558 4639
rect 15575 4622 15581 4639
rect 15552 4614 15581 4622
rect 15596 4809 15625 4814
rect 15596 4792 15602 4809
rect 15619 4792 15625 4809
rect 15596 4775 15625 4792
rect 15596 4758 15602 4775
rect 15619 4758 15625 4775
rect 15596 4741 15625 4758
rect 15596 4724 15602 4741
rect 15619 4724 15625 4741
rect 15596 4707 15625 4724
rect 15596 4690 15602 4707
rect 15619 4690 15625 4707
rect 15596 4673 15625 4690
rect 15596 4656 15602 4673
rect 15619 4656 15625 4673
rect 15596 4639 15625 4656
rect 15596 4622 15602 4639
rect 15619 4622 15625 4639
rect 15596 4614 15625 4622
rect 15640 4809 15669 4814
rect 15640 4792 15646 4809
rect 15663 4792 15669 4809
rect 15640 4775 15669 4792
rect 15640 4758 15646 4775
rect 15663 4758 15669 4775
rect 15640 4741 15669 4758
rect 15640 4724 15646 4741
rect 15663 4724 15669 4741
rect 15640 4707 15669 4724
rect 15640 4690 15646 4707
rect 15663 4690 15669 4707
rect 15640 4673 15669 4690
rect 15640 4656 15646 4673
rect 15663 4656 15669 4673
rect 15640 4639 15669 4656
rect 15640 4622 15646 4639
rect 15663 4622 15669 4639
rect 15640 4614 15669 4622
<< ndiffc >>
rect 13067 7646 13084 7663
rect 13067 7612 13084 7629
rect 13067 7578 13084 7595
rect 13147 7646 13164 7663
rect 13147 7612 13164 7629
rect 13147 7578 13164 7595
rect 13191 7646 13208 7663
rect 13191 7612 13208 7629
rect 13191 7578 13208 7595
rect 13235 7646 13252 7663
rect 13235 7612 13252 7629
rect 13235 7578 13252 7595
rect 13315 7646 13332 7663
rect 13315 7612 13332 7629
rect 13315 7578 13332 7595
rect 13678 7646 13695 7663
rect 13678 7612 13695 7629
rect 13678 7578 13695 7595
rect 13758 7646 13775 7663
rect 13758 7612 13775 7629
rect 13758 7578 13775 7595
rect 13802 7646 13819 7663
rect 13802 7612 13819 7629
rect 13802 7578 13819 7595
rect 13846 7646 13863 7663
rect 13846 7612 13863 7629
rect 13846 7578 13863 7595
rect 13926 7646 13943 7663
rect 13926 7612 13943 7629
rect 13926 7578 13943 7595
rect 14256 7646 14273 7663
rect 14256 7612 14273 7629
rect 14256 7578 14273 7595
rect 14336 7646 14353 7663
rect 14336 7612 14353 7629
rect 14336 7578 14353 7595
rect 14380 7646 14397 7663
rect 14380 7612 14397 7629
rect 14380 7578 14397 7595
rect 14424 7646 14441 7663
rect 14424 7612 14441 7629
rect 14424 7578 14441 7595
rect 14504 7646 14521 7663
rect 14504 7612 14521 7629
rect 14504 7578 14521 7595
rect 14867 7646 14884 7663
rect 14867 7612 14884 7629
rect 14867 7578 14884 7595
rect 14947 7646 14964 7663
rect 14947 7612 14964 7629
rect 14947 7578 14964 7595
rect 14991 7646 15008 7663
rect 14991 7612 15008 7629
rect 14991 7578 15008 7595
rect 15035 7646 15052 7663
rect 15035 7612 15052 7629
rect 15035 7578 15052 7595
rect 15115 7646 15132 7663
rect 15115 7612 15132 7629
rect 15115 7578 15132 7595
rect 15478 7646 15495 7663
rect 15478 7612 15495 7629
rect 15478 7578 15495 7595
rect 15558 7646 15575 7663
rect 15558 7612 15575 7629
rect 15558 7578 15575 7595
rect 15602 7646 15619 7663
rect 15602 7612 15619 7629
rect 15602 7578 15619 7595
rect 15646 7646 15663 7663
rect 15646 7612 15663 7629
rect 15646 7578 15663 7595
rect 15726 7646 15743 7663
rect 15726 7612 15743 7629
rect 15726 7578 15743 7595
rect 12456 6996 12473 7013
rect 12456 6962 12473 6979
rect 12456 6928 12473 6945
rect 12536 6996 12553 7013
rect 12536 6962 12553 6979
rect 12536 6928 12553 6945
rect 12580 6996 12597 7013
rect 12580 6962 12597 6979
rect 12580 6928 12597 6945
rect 12624 6996 12641 7013
rect 12624 6962 12641 6979
rect 12624 6928 12641 6945
rect 12704 6996 12721 7013
rect 12704 6962 12721 6979
rect 12704 6928 12721 6945
rect 13067 6996 13084 7013
rect 13067 6962 13084 6979
rect 13067 6928 13084 6945
rect 13147 6996 13164 7013
rect 13147 6962 13164 6979
rect 13147 6928 13164 6945
rect 13191 6996 13208 7013
rect 13191 6962 13208 6979
rect 13191 6928 13208 6945
rect 13235 6996 13252 7013
rect 13235 6962 13252 6979
rect 13235 6928 13252 6945
rect 13315 6996 13332 7013
rect 13315 6962 13332 6979
rect 13315 6928 13332 6945
rect 13678 6996 13695 7013
rect 13678 6962 13695 6979
rect 13678 6928 13695 6945
rect 13758 6996 13775 7013
rect 13758 6962 13775 6979
rect 13758 6928 13775 6945
rect 13802 6996 13819 7013
rect 13802 6962 13819 6979
rect 13802 6928 13819 6945
rect 13846 6996 13863 7013
rect 13846 6962 13863 6979
rect 13846 6928 13863 6945
rect 13926 6996 13943 7013
rect 13926 6962 13943 6979
rect 13926 6928 13943 6945
rect 14256 6996 14273 7013
rect 14256 6962 14273 6979
rect 14256 6928 14273 6945
rect 14336 6996 14353 7013
rect 14336 6962 14353 6979
rect 14336 6928 14353 6945
rect 14380 6996 14397 7013
rect 14380 6962 14397 6979
rect 14380 6928 14397 6945
rect 14424 6996 14441 7013
rect 14424 6962 14441 6979
rect 14424 6928 14441 6945
rect 14504 6996 14521 7013
rect 14504 6962 14521 6979
rect 14504 6928 14521 6945
rect 14867 6996 14884 7013
rect 14867 6962 14884 6979
rect 14867 6928 14884 6945
rect 14947 6996 14964 7013
rect 14947 6962 14964 6979
rect 14947 6928 14964 6945
rect 14991 6996 15008 7013
rect 14991 6962 15008 6979
rect 14991 6928 15008 6945
rect 15035 6996 15052 7013
rect 15035 6962 15052 6979
rect 15035 6928 15052 6945
rect 15115 6996 15132 7013
rect 15115 6962 15132 6979
rect 15115 6928 15132 6945
rect 15478 6996 15495 7013
rect 15478 6962 15495 6979
rect 15478 6928 15495 6945
rect 15558 6996 15575 7013
rect 15558 6962 15575 6979
rect 15558 6928 15575 6945
rect 15602 6996 15619 7013
rect 15602 6962 15619 6979
rect 15602 6928 15619 6945
rect 15646 6996 15663 7013
rect 15646 6962 15663 6979
rect 15646 6928 15663 6945
rect 15726 6996 15743 7013
rect 15726 6962 15743 6979
rect 15726 6928 15743 6945
rect 12456 6356 12473 6373
rect 12456 6322 12473 6339
rect 12456 6288 12473 6305
rect 12536 6356 12553 6373
rect 12536 6322 12553 6339
rect 12536 6288 12553 6305
rect 12580 6356 12597 6373
rect 12580 6322 12597 6339
rect 12580 6288 12597 6305
rect 12624 6356 12641 6373
rect 12624 6322 12641 6339
rect 12624 6288 12641 6305
rect 12704 6356 12721 6373
rect 12704 6322 12721 6339
rect 12704 6288 12721 6305
rect 13067 6356 13084 6373
rect 13067 6322 13084 6339
rect 13067 6288 13084 6305
rect 13147 6356 13164 6373
rect 13147 6322 13164 6339
rect 13147 6288 13164 6305
rect 13191 6356 13208 6373
rect 13191 6322 13208 6339
rect 13191 6288 13208 6305
rect 13235 6356 13252 6373
rect 13235 6322 13252 6339
rect 13235 6288 13252 6305
rect 13315 6356 13332 6373
rect 13315 6322 13332 6339
rect 13315 6288 13332 6305
rect 13678 6356 13695 6373
rect 13678 6322 13695 6339
rect 13678 6288 13695 6305
rect 13758 6356 13775 6373
rect 13758 6322 13775 6339
rect 13758 6288 13775 6305
rect 13802 6356 13819 6373
rect 13802 6322 13819 6339
rect 13802 6288 13819 6305
rect 13846 6356 13863 6373
rect 13846 6322 13863 6339
rect 13846 6288 13863 6305
rect 13926 6356 13943 6373
rect 13926 6322 13943 6339
rect 13926 6288 13943 6305
rect 14256 6356 14273 6373
rect 14256 6322 14273 6339
rect 14256 6288 14273 6305
rect 14336 6356 14353 6373
rect 14336 6322 14353 6339
rect 14336 6288 14353 6305
rect 14380 6356 14397 6373
rect 14380 6322 14397 6339
rect 14380 6288 14397 6305
rect 14424 6356 14441 6373
rect 14424 6322 14441 6339
rect 14424 6288 14441 6305
rect 14504 6356 14521 6373
rect 14504 6322 14521 6339
rect 14504 6288 14521 6305
rect 14867 6356 14884 6373
rect 14867 6322 14884 6339
rect 14867 6288 14884 6305
rect 14947 6356 14964 6373
rect 14947 6322 14964 6339
rect 14947 6288 14964 6305
rect 14991 6356 15008 6373
rect 14991 6322 15008 6339
rect 14991 6288 15008 6305
rect 15035 6356 15052 6373
rect 15035 6322 15052 6339
rect 15035 6288 15052 6305
rect 15115 6356 15132 6373
rect 15115 6322 15132 6339
rect 15115 6288 15132 6305
rect 15478 6356 15495 6373
rect 15478 6322 15495 6339
rect 15478 6288 15495 6305
rect 15558 6356 15575 6373
rect 15558 6322 15575 6339
rect 15558 6288 15575 6305
rect 15602 6356 15619 6373
rect 15602 6322 15619 6339
rect 15602 6288 15619 6305
rect 15646 6356 15663 6373
rect 15646 6322 15663 6339
rect 15646 6288 15663 6305
rect 15726 6356 15743 6373
rect 15726 6322 15743 6339
rect 15726 6288 15743 6305
rect 12456 5706 12473 5723
rect 12456 5672 12473 5689
rect 12456 5638 12473 5655
rect 12536 5706 12553 5723
rect 12536 5672 12553 5689
rect 12536 5638 12553 5655
rect 12580 5706 12597 5723
rect 12580 5672 12597 5689
rect 12580 5638 12597 5655
rect 12624 5706 12641 5723
rect 12624 5672 12641 5689
rect 12624 5638 12641 5655
rect 12704 5706 12721 5723
rect 12704 5672 12721 5689
rect 12704 5638 12721 5655
rect 13067 5706 13084 5723
rect 13067 5672 13084 5689
rect 13067 5638 13084 5655
rect 13147 5706 13164 5723
rect 13147 5672 13164 5689
rect 13147 5638 13164 5655
rect 13191 5706 13208 5723
rect 13191 5672 13208 5689
rect 13191 5638 13208 5655
rect 13235 5706 13252 5723
rect 13235 5672 13252 5689
rect 13235 5638 13252 5655
rect 13315 5706 13332 5723
rect 13315 5672 13332 5689
rect 13315 5638 13332 5655
rect 13678 5706 13695 5723
rect 13678 5672 13695 5689
rect 13678 5638 13695 5655
rect 13758 5706 13775 5723
rect 13758 5672 13775 5689
rect 13758 5638 13775 5655
rect 13802 5706 13819 5723
rect 13802 5672 13819 5689
rect 13802 5638 13819 5655
rect 13846 5706 13863 5723
rect 13846 5672 13863 5689
rect 13846 5638 13863 5655
rect 13926 5706 13943 5723
rect 13926 5672 13943 5689
rect 13926 5638 13943 5655
rect 14256 5706 14273 5723
rect 14256 5672 14273 5689
rect 14256 5638 14273 5655
rect 14336 5706 14353 5723
rect 14336 5672 14353 5689
rect 14336 5638 14353 5655
rect 14380 5706 14397 5723
rect 14380 5672 14397 5689
rect 14380 5638 14397 5655
rect 14424 5706 14441 5723
rect 14424 5672 14441 5689
rect 14424 5638 14441 5655
rect 14504 5706 14521 5723
rect 14504 5672 14521 5689
rect 14504 5638 14521 5655
rect 14867 5706 14884 5723
rect 14867 5672 14884 5689
rect 14867 5638 14884 5655
rect 14947 5706 14964 5723
rect 14947 5672 14964 5689
rect 14947 5638 14964 5655
rect 14991 5706 15008 5723
rect 14991 5672 15008 5689
rect 14991 5638 15008 5655
rect 15035 5706 15052 5723
rect 15035 5672 15052 5689
rect 15035 5638 15052 5655
rect 15115 5706 15132 5723
rect 15115 5672 15132 5689
rect 15115 5638 15132 5655
rect 15478 5706 15495 5723
rect 15478 5672 15495 5689
rect 15478 5638 15495 5655
rect 15558 5706 15575 5723
rect 15558 5672 15575 5689
rect 15558 5638 15575 5655
rect 15602 5706 15619 5723
rect 15602 5672 15619 5689
rect 15602 5638 15619 5655
rect 15646 5706 15663 5723
rect 15646 5672 15663 5689
rect 15646 5638 15663 5655
rect 15726 5706 15743 5723
rect 15726 5672 15743 5689
rect 15726 5638 15743 5655
rect 12456 5056 12473 5073
rect 12456 5022 12473 5039
rect 12456 4988 12473 5005
rect 12536 5056 12553 5073
rect 12536 5022 12553 5039
rect 12536 4988 12553 5005
rect 12580 5056 12597 5073
rect 12580 5022 12597 5039
rect 12580 4988 12597 5005
rect 12624 5056 12641 5073
rect 12624 5022 12641 5039
rect 12624 4988 12641 5005
rect 12704 5056 12721 5073
rect 12704 5022 12721 5039
rect 12704 4988 12721 5005
rect 13067 5056 13084 5073
rect 13067 5022 13084 5039
rect 13067 4988 13084 5005
rect 13147 5056 13164 5073
rect 13147 5022 13164 5039
rect 13147 4988 13164 5005
rect 13191 5056 13208 5073
rect 13191 5022 13208 5039
rect 13191 4988 13208 5005
rect 13235 5056 13252 5073
rect 13235 5022 13252 5039
rect 13235 4988 13252 5005
rect 13315 5056 13332 5073
rect 13315 5022 13332 5039
rect 13315 4988 13332 5005
rect 13678 5056 13695 5073
rect 13678 5022 13695 5039
rect 13678 4988 13695 5005
rect 13758 5056 13775 5073
rect 13758 5022 13775 5039
rect 13758 4988 13775 5005
rect 13802 5056 13819 5073
rect 13802 5022 13819 5039
rect 13802 4988 13819 5005
rect 13846 5056 13863 5073
rect 13846 5022 13863 5039
rect 13846 4988 13863 5005
rect 13926 5056 13943 5073
rect 13926 5022 13943 5039
rect 13926 4988 13943 5005
rect 14256 5056 14273 5073
rect 14256 5022 14273 5039
rect 14256 4988 14273 5005
rect 14336 5056 14353 5073
rect 14336 5022 14353 5039
rect 14336 4988 14353 5005
rect 14380 5056 14397 5073
rect 14380 5022 14397 5039
rect 14380 4988 14397 5005
rect 14424 5056 14441 5073
rect 14424 5022 14441 5039
rect 14424 4988 14441 5005
rect 14504 5056 14521 5073
rect 14504 5022 14521 5039
rect 14504 4988 14521 5005
rect 14867 5056 14884 5073
rect 14867 5022 14884 5039
rect 14867 4988 14884 5005
rect 14947 5056 14964 5073
rect 14947 5022 14964 5039
rect 14947 4988 14964 5005
rect 14991 5056 15008 5073
rect 14991 5022 15008 5039
rect 14991 4988 15008 5005
rect 15035 5056 15052 5073
rect 15035 5022 15052 5039
rect 15035 4988 15052 5005
rect 15115 5056 15132 5073
rect 15115 5022 15132 5039
rect 15115 4988 15132 5005
rect 15478 5056 15495 5073
rect 15478 5022 15495 5039
rect 15478 4988 15495 5005
rect 15558 5056 15575 5073
rect 15558 5022 15575 5039
rect 15558 4988 15575 5005
rect 15602 5056 15619 5073
rect 15602 5022 15619 5039
rect 15602 4988 15619 5005
rect 15646 5056 15663 5073
rect 15646 5022 15663 5039
rect 15646 4988 15663 5005
rect 15726 5056 15743 5073
rect 15726 5022 15743 5039
rect 15726 4988 15743 5005
rect 12456 4416 12473 4433
rect 12456 4382 12473 4399
rect 12456 4348 12473 4365
rect 12536 4416 12553 4433
rect 12536 4382 12553 4399
rect 12536 4348 12553 4365
rect 12580 4416 12597 4433
rect 12580 4382 12597 4399
rect 12580 4348 12597 4365
rect 12624 4416 12641 4433
rect 12624 4382 12641 4399
rect 12624 4348 12641 4365
rect 12704 4416 12721 4433
rect 12704 4382 12721 4399
rect 12704 4348 12721 4365
rect 13067 4416 13084 4433
rect 13067 4382 13084 4399
rect 13067 4348 13084 4365
rect 13147 4416 13164 4433
rect 13147 4382 13164 4399
rect 13147 4348 13164 4365
rect 13191 4416 13208 4433
rect 13191 4382 13208 4399
rect 13191 4348 13208 4365
rect 13235 4416 13252 4433
rect 13235 4382 13252 4399
rect 13235 4348 13252 4365
rect 13315 4416 13332 4433
rect 13315 4382 13332 4399
rect 13315 4348 13332 4365
rect 13678 4416 13695 4433
rect 13678 4382 13695 4399
rect 13678 4348 13695 4365
rect 13758 4416 13775 4433
rect 13758 4382 13775 4399
rect 13758 4348 13775 4365
rect 13802 4416 13819 4433
rect 13802 4382 13819 4399
rect 13802 4348 13819 4365
rect 13846 4416 13863 4433
rect 13846 4382 13863 4399
rect 13846 4348 13863 4365
rect 13926 4416 13943 4433
rect 13926 4382 13943 4399
rect 13926 4348 13943 4365
rect 14256 4416 14273 4433
rect 14256 4382 14273 4399
rect 14256 4348 14273 4365
rect 14336 4416 14353 4433
rect 14336 4382 14353 4399
rect 14336 4348 14353 4365
rect 14380 4416 14397 4433
rect 14380 4382 14397 4399
rect 14380 4348 14397 4365
rect 14424 4416 14441 4433
rect 14424 4382 14441 4399
rect 14424 4348 14441 4365
rect 14504 4416 14521 4433
rect 14504 4382 14521 4399
rect 14504 4348 14521 4365
rect 14867 4416 14884 4433
rect 14867 4382 14884 4399
rect 14867 4348 14884 4365
rect 14947 4416 14964 4433
rect 14947 4382 14964 4399
rect 14947 4348 14964 4365
rect 14991 4416 15008 4433
rect 14991 4382 15008 4399
rect 14991 4348 15008 4365
rect 15035 4416 15052 4433
rect 15035 4382 15052 4399
rect 15035 4348 15052 4365
rect 15115 4416 15132 4433
rect 15115 4382 15132 4399
rect 15115 4348 15132 4365
rect 15478 4416 15495 4433
rect 15478 4382 15495 4399
rect 15478 4348 15495 4365
rect 15558 4416 15575 4433
rect 15558 4382 15575 4399
rect 15558 4348 15575 4365
rect 15602 4416 15619 4433
rect 15602 4382 15619 4399
rect 15602 4348 15619 4365
rect 15646 4416 15663 4433
rect 15646 4382 15663 4399
rect 15646 4348 15663 4365
rect 15726 4416 15743 4433
rect 15726 4382 15743 4399
rect 15726 4348 15743 4365
<< pdiffc >>
rect 13147 8022 13164 8039
rect 13147 7988 13164 8005
rect 13147 7954 13164 7971
rect 13147 7920 13164 7937
rect 13147 7886 13164 7903
rect 13147 7852 13164 7869
rect 13191 8022 13208 8039
rect 13191 7988 13208 8005
rect 13191 7954 13208 7971
rect 13191 7920 13208 7937
rect 13191 7886 13208 7903
rect 13191 7852 13208 7869
rect 13235 8022 13252 8039
rect 13235 7988 13252 8005
rect 13235 7954 13252 7971
rect 13235 7920 13252 7937
rect 13235 7886 13252 7903
rect 13235 7852 13252 7869
rect 13758 8022 13775 8039
rect 13758 7988 13775 8005
rect 13758 7954 13775 7971
rect 13758 7920 13775 7937
rect 13758 7886 13775 7903
rect 13758 7852 13775 7869
rect 13802 8022 13819 8039
rect 13802 7988 13819 8005
rect 13802 7954 13819 7971
rect 13802 7920 13819 7937
rect 13802 7886 13819 7903
rect 13802 7852 13819 7869
rect 13846 8022 13863 8039
rect 13846 7988 13863 8005
rect 13846 7954 13863 7971
rect 13846 7920 13863 7937
rect 13846 7886 13863 7903
rect 13846 7852 13863 7869
rect 14336 8022 14353 8039
rect 14336 7988 14353 8005
rect 14336 7954 14353 7971
rect 14336 7920 14353 7937
rect 14336 7886 14353 7903
rect 14336 7852 14353 7869
rect 14380 8022 14397 8039
rect 14380 7988 14397 8005
rect 14380 7954 14397 7971
rect 14380 7920 14397 7937
rect 14380 7886 14397 7903
rect 14380 7852 14397 7869
rect 14424 8022 14441 8039
rect 14424 7988 14441 8005
rect 14424 7954 14441 7971
rect 14424 7920 14441 7937
rect 14424 7886 14441 7903
rect 14424 7852 14441 7869
rect 14947 8022 14964 8039
rect 14947 7988 14964 8005
rect 14947 7954 14964 7971
rect 14947 7920 14964 7937
rect 14947 7886 14964 7903
rect 14947 7852 14964 7869
rect 14991 8022 15008 8039
rect 14991 7988 15008 8005
rect 14991 7954 15008 7971
rect 14991 7920 15008 7937
rect 14991 7886 15008 7903
rect 14991 7852 15008 7869
rect 15035 8022 15052 8039
rect 15035 7988 15052 8005
rect 15035 7954 15052 7971
rect 15035 7920 15052 7937
rect 15035 7886 15052 7903
rect 15035 7852 15052 7869
rect 15558 8022 15575 8039
rect 15558 7988 15575 8005
rect 15558 7954 15575 7971
rect 15558 7920 15575 7937
rect 15558 7886 15575 7903
rect 15558 7852 15575 7869
rect 15602 8022 15619 8039
rect 15602 7988 15619 8005
rect 15602 7954 15619 7971
rect 15602 7920 15619 7937
rect 15602 7886 15619 7903
rect 15602 7852 15619 7869
rect 15646 8022 15663 8039
rect 15646 7988 15663 8005
rect 15646 7954 15663 7971
rect 15646 7920 15663 7937
rect 15646 7886 15663 7903
rect 15646 7852 15663 7869
rect 12536 7372 12553 7389
rect 12536 7338 12553 7355
rect 12536 7304 12553 7321
rect 12536 7270 12553 7287
rect 12536 7236 12553 7253
rect 12536 7202 12553 7219
rect 12580 7372 12597 7389
rect 12580 7338 12597 7355
rect 12580 7304 12597 7321
rect 12580 7270 12597 7287
rect 12580 7236 12597 7253
rect 12580 7202 12597 7219
rect 12624 7372 12641 7389
rect 12624 7338 12641 7355
rect 12624 7304 12641 7321
rect 12624 7270 12641 7287
rect 12624 7236 12641 7253
rect 12624 7202 12641 7219
rect 13147 7372 13164 7389
rect 13147 7338 13164 7355
rect 13147 7304 13164 7321
rect 13147 7270 13164 7287
rect 13147 7236 13164 7253
rect 13147 7202 13164 7219
rect 13191 7372 13208 7389
rect 13191 7338 13208 7355
rect 13191 7304 13208 7321
rect 13191 7270 13208 7287
rect 13191 7236 13208 7253
rect 13191 7202 13208 7219
rect 13235 7372 13252 7389
rect 13235 7338 13252 7355
rect 13235 7304 13252 7321
rect 13235 7270 13252 7287
rect 13235 7236 13252 7253
rect 13235 7202 13252 7219
rect 13758 7372 13775 7389
rect 13758 7338 13775 7355
rect 13758 7304 13775 7321
rect 13758 7270 13775 7287
rect 13758 7236 13775 7253
rect 13758 7202 13775 7219
rect 13802 7372 13819 7389
rect 13802 7338 13819 7355
rect 13802 7304 13819 7321
rect 13802 7270 13819 7287
rect 13802 7236 13819 7253
rect 13802 7202 13819 7219
rect 13846 7372 13863 7389
rect 13846 7338 13863 7355
rect 13846 7304 13863 7321
rect 13846 7270 13863 7287
rect 13846 7236 13863 7253
rect 13846 7202 13863 7219
rect 14336 7372 14353 7389
rect 14336 7338 14353 7355
rect 14336 7304 14353 7321
rect 14336 7270 14353 7287
rect 14336 7236 14353 7253
rect 14336 7202 14353 7219
rect 14380 7372 14397 7389
rect 14380 7338 14397 7355
rect 14380 7304 14397 7321
rect 14380 7270 14397 7287
rect 14380 7236 14397 7253
rect 14380 7202 14397 7219
rect 14424 7372 14441 7389
rect 14424 7338 14441 7355
rect 14424 7304 14441 7321
rect 14424 7270 14441 7287
rect 14424 7236 14441 7253
rect 14424 7202 14441 7219
rect 14947 7372 14964 7389
rect 14947 7338 14964 7355
rect 14947 7304 14964 7321
rect 14947 7270 14964 7287
rect 14947 7236 14964 7253
rect 14947 7202 14964 7219
rect 14991 7372 15008 7389
rect 14991 7338 15008 7355
rect 14991 7304 15008 7321
rect 14991 7270 15008 7287
rect 14991 7236 15008 7253
rect 14991 7202 15008 7219
rect 15035 7372 15052 7389
rect 15035 7338 15052 7355
rect 15035 7304 15052 7321
rect 15035 7270 15052 7287
rect 15035 7236 15052 7253
rect 15035 7202 15052 7219
rect 15558 7372 15575 7389
rect 15558 7338 15575 7355
rect 15558 7304 15575 7321
rect 15558 7270 15575 7287
rect 15558 7236 15575 7253
rect 15558 7202 15575 7219
rect 15602 7372 15619 7389
rect 15602 7338 15619 7355
rect 15602 7304 15619 7321
rect 15602 7270 15619 7287
rect 15602 7236 15619 7253
rect 15602 7202 15619 7219
rect 15646 7372 15663 7389
rect 15646 7338 15663 7355
rect 15646 7304 15663 7321
rect 15646 7270 15663 7287
rect 15646 7236 15663 7253
rect 15646 7202 15663 7219
rect 12536 6732 12553 6749
rect 12536 6698 12553 6715
rect 12536 6664 12553 6681
rect 12536 6630 12553 6647
rect 12536 6596 12553 6613
rect 12536 6562 12553 6579
rect 12580 6732 12597 6749
rect 12580 6698 12597 6715
rect 12580 6664 12597 6681
rect 12580 6630 12597 6647
rect 12580 6596 12597 6613
rect 12580 6562 12597 6579
rect 12624 6732 12641 6749
rect 12624 6698 12641 6715
rect 12624 6664 12641 6681
rect 12624 6630 12641 6647
rect 12624 6596 12641 6613
rect 12624 6562 12641 6579
rect 13147 6732 13164 6749
rect 13147 6698 13164 6715
rect 13147 6664 13164 6681
rect 13147 6630 13164 6647
rect 13147 6596 13164 6613
rect 13147 6562 13164 6579
rect 13191 6732 13208 6749
rect 13191 6698 13208 6715
rect 13191 6664 13208 6681
rect 13191 6630 13208 6647
rect 13191 6596 13208 6613
rect 13191 6562 13208 6579
rect 13235 6732 13252 6749
rect 13235 6698 13252 6715
rect 13235 6664 13252 6681
rect 13235 6630 13252 6647
rect 13235 6596 13252 6613
rect 13235 6562 13252 6579
rect 13758 6732 13775 6749
rect 13758 6698 13775 6715
rect 13758 6664 13775 6681
rect 13758 6630 13775 6647
rect 13758 6596 13775 6613
rect 13758 6562 13775 6579
rect 13802 6732 13819 6749
rect 13802 6698 13819 6715
rect 13802 6664 13819 6681
rect 13802 6630 13819 6647
rect 13802 6596 13819 6613
rect 13802 6562 13819 6579
rect 13846 6732 13863 6749
rect 13846 6698 13863 6715
rect 13846 6664 13863 6681
rect 13846 6630 13863 6647
rect 13846 6596 13863 6613
rect 13846 6562 13863 6579
rect 14336 6732 14353 6749
rect 14336 6698 14353 6715
rect 14336 6664 14353 6681
rect 14336 6630 14353 6647
rect 14336 6596 14353 6613
rect 14336 6562 14353 6579
rect 14380 6732 14397 6749
rect 14380 6698 14397 6715
rect 14380 6664 14397 6681
rect 14380 6630 14397 6647
rect 14380 6596 14397 6613
rect 14380 6562 14397 6579
rect 14424 6732 14441 6749
rect 14424 6698 14441 6715
rect 14424 6664 14441 6681
rect 14424 6630 14441 6647
rect 14424 6596 14441 6613
rect 14424 6562 14441 6579
rect 14947 6732 14964 6749
rect 14947 6698 14964 6715
rect 14947 6664 14964 6681
rect 14947 6630 14964 6647
rect 14947 6596 14964 6613
rect 14947 6562 14964 6579
rect 14991 6732 15008 6749
rect 14991 6698 15008 6715
rect 14991 6664 15008 6681
rect 14991 6630 15008 6647
rect 14991 6596 15008 6613
rect 14991 6562 15008 6579
rect 15035 6732 15052 6749
rect 15035 6698 15052 6715
rect 15035 6664 15052 6681
rect 15035 6630 15052 6647
rect 15035 6596 15052 6613
rect 15035 6562 15052 6579
rect 15558 6732 15575 6749
rect 15558 6698 15575 6715
rect 15558 6664 15575 6681
rect 15558 6630 15575 6647
rect 15558 6596 15575 6613
rect 15558 6562 15575 6579
rect 15602 6732 15619 6749
rect 15602 6698 15619 6715
rect 15602 6664 15619 6681
rect 15602 6630 15619 6647
rect 15602 6596 15619 6613
rect 15602 6562 15619 6579
rect 15646 6732 15663 6749
rect 15646 6698 15663 6715
rect 15646 6664 15663 6681
rect 15646 6630 15663 6647
rect 15646 6596 15663 6613
rect 15646 6562 15663 6579
rect 12536 6082 12553 6099
rect 12536 6048 12553 6065
rect 12536 6014 12553 6031
rect 12536 5980 12553 5997
rect 12536 5946 12553 5963
rect 12536 5912 12553 5929
rect 12580 6082 12597 6099
rect 12580 6048 12597 6065
rect 12580 6014 12597 6031
rect 12580 5980 12597 5997
rect 12580 5946 12597 5963
rect 12580 5912 12597 5929
rect 12624 6082 12641 6099
rect 12624 6048 12641 6065
rect 12624 6014 12641 6031
rect 12624 5980 12641 5997
rect 12624 5946 12641 5963
rect 12624 5912 12641 5929
rect 13147 6082 13164 6099
rect 13147 6048 13164 6065
rect 13147 6014 13164 6031
rect 13147 5980 13164 5997
rect 13147 5946 13164 5963
rect 13147 5912 13164 5929
rect 13191 6082 13208 6099
rect 13191 6048 13208 6065
rect 13191 6014 13208 6031
rect 13191 5980 13208 5997
rect 13191 5946 13208 5963
rect 13191 5912 13208 5929
rect 13235 6082 13252 6099
rect 13235 6048 13252 6065
rect 13235 6014 13252 6031
rect 13235 5980 13252 5997
rect 13235 5946 13252 5963
rect 13235 5912 13252 5929
rect 13758 6082 13775 6099
rect 13758 6048 13775 6065
rect 13758 6014 13775 6031
rect 13758 5980 13775 5997
rect 13758 5946 13775 5963
rect 13758 5912 13775 5929
rect 13802 6082 13819 6099
rect 13802 6048 13819 6065
rect 13802 6014 13819 6031
rect 13802 5980 13819 5997
rect 13802 5946 13819 5963
rect 13802 5912 13819 5929
rect 13846 6082 13863 6099
rect 13846 6048 13863 6065
rect 13846 6014 13863 6031
rect 13846 5980 13863 5997
rect 13846 5946 13863 5963
rect 13846 5912 13863 5929
rect 14336 6082 14353 6099
rect 14336 6048 14353 6065
rect 14336 6014 14353 6031
rect 14336 5980 14353 5997
rect 14336 5946 14353 5963
rect 14336 5912 14353 5929
rect 14380 6082 14397 6099
rect 14380 6048 14397 6065
rect 14380 6014 14397 6031
rect 14380 5980 14397 5997
rect 14380 5946 14397 5963
rect 14380 5912 14397 5929
rect 14424 6082 14441 6099
rect 14424 6048 14441 6065
rect 14424 6014 14441 6031
rect 14424 5980 14441 5997
rect 14424 5946 14441 5963
rect 14424 5912 14441 5929
rect 14947 6082 14964 6099
rect 14947 6048 14964 6065
rect 14947 6014 14964 6031
rect 14947 5980 14964 5997
rect 14947 5946 14964 5963
rect 14947 5912 14964 5929
rect 14991 6082 15008 6099
rect 14991 6048 15008 6065
rect 14991 6014 15008 6031
rect 14991 5980 15008 5997
rect 14991 5946 15008 5963
rect 14991 5912 15008 5929
rect 15035 6082 15052 6099
rect 15035 6048 15052 6065
rect 15035 6014 15052 6031
rect 15035 5980 15052 5997
rect 15035 5946 15052 5963
rect 15035 5912 15052 5929
rect 15558 6082 15575 6099
rect 15558 6048 15575 6065
rect 15558 6014 15575 6031
rect 15558 5980 15575 5997
rect 15558 5946 15575 5963
rect 15558 5912 15575 5929
rect 15602 6082 15619 6099
rect 15602 6048 15619 6065
rect 15602 6014 15619 6031
rect 15602 5980 15619 5997
rect 15602 5946 15619 5963
rect 15602 5912 15619 5929
rect 15646 6082 15663 6099
rect 15646 6048 15663 6065
rect 15646 6014 15663 6031
rect 15646 5980 15663 5997
rect 15646 5946 15663 5963
rect 15646 5912 15663 5929
rect 12536 5432 12553 5449
rect 12536 5398 12553 5415
rect 12536 5364 12553 5381
rect 12536 5330 12553 5347
rect 12536 5296 12553 5313
rect 12536 5262 12553 5279
rect 12580 5432 12597 5449
rect 12580 5398 12597 5415
rect 12580 5364 12597 5381
rect 12580 5330 12597 5347
rect 12580 5296 12597 5313
rect 12580 5262 12597 5279
rect 12624 5432 12641 5449
rect 12624 5398 12641 5415
rect 12624 5364 12641 5381
rect 12624 5330 12641 5347
rect 12624 5296 12641 5313
rect 12624 5262 12641 5279
rect 13147 5432 13164 5449
rect 13147 5398 13164 5415
rect 13147 5364 13164 5381
rect 13147 5330 13164 5347
rect 13147 5296 13164 5313
rect 13147 5262 13164 5279
rect 13191 5432 13208 5449
rect 13191 5398 13208 5415
rect 13191 5364 13208 5381
rect 13191 5330 13208 5347
rect 13191 5296 13208 5313
rect 13191 5262 13208 5279
rect 13235 5432 13252 5449
rect 13235 5398 13252 5415
rect 13235 5364 13252 5381
rect 13235 5330 13252 5347
rect 13235 5296 13252 5313
rect 13235 5262 13252 5279
rect 13758 5432 13775 5449
rect 13758 5398 13775 5415
rect 13758 5364 13775 5381
rect 13758 5330 13775 5347
rect 13758 5296 13775 5313
rect 13758 5262 13775 5279
rect 13802 5432 13819 5449
rect 13802 5398 13819 5415
rect 13802 5364 13819 5381
rect 13802 5330 13819 5347
rect 13802 5296 13819 5313
rect 13802 5262 13819 5279
rect 13846 5432 13863 5449
rect 13846 5398 13863 5415
rect 13846 5364 13863 5381
rect 13846 5330 13863 5347
rect 13846 5296 13863 5313
rect 13846 5262 13863 5279
rect 14336 5432 14353 5449
rect 14336 5398 14353 5415
rect 14336 5364 14353 5381
rect 14336 5330 14353 5347
rect 14336 5296 14353 5313
rect 14336 5262 14353 5279
rect 14380 5432 14397 5449
rect 14380 5398 14397 5415
rect 14380 5364 14397 5381
rect 14380 5330 14397 5347
rect 14380 5296 14397 5313
rect 14380 5262 14397 5279
rect 14424 5432 14441 5449
rect 14424 5398 14441 5415
rect 14424 5364 14441 5381
rect 14424 5330 14441 5347
rect 14424 5296 14441 5313
rect 14424 5262 14441 5279
rect 14947 5432 14964 5449
rect 14947 5398 14964 5415
rect 14947 5364 14964 5381
rect 14947 5330 14964 5347
rect 14947 5296 14964 5313
rect 14947 5262 14964 5279
rect 14991 5432 15008 5449
rect 14991 5398 15008 5415
rect 14991 5364 15008 5381
rect 14991 5330 15008 5347
rect 14991 5296 15008 5313
rect 14991 5262 15008 5279
rect 15035 5432 15052 5449
rect 15035 5398 15052 5415
rect 15035 5364 15052 5381
rect 15035 5330 15052 5347
rect 15035 5296 15052 5313
rect 15035 5262 15052 5279
rect 15558 5432 15575 5449
rect 15558 5398 15575 5415
rect 15558 5364 15575 5381
rect 15558 5330 15575 5347
rect 15558 5296 15575 5313
rect 15558 5262 15575 5279
rect 15602 5432 15619 5449
rect 15602 5398 15619 5415
rect 15602 5364 15619 5381
rect 15602 5330 15619 5347
rect 15602 5296 15619 5313
rect 15602 5262 15619 5279
rect 15646 5432 15663 5449
rect 15646 5398 15663 5415
rect 15646 5364 15663 5381
rect 15646 5330 15663 5347
rect 15646 5296 15663 5313
rect 15646 5262 15663 5279
rect 12536 4792 12553 4809
rect 12536 4758 12553 4775
rect 12536 4724 12553 4741
rect 12536 4690 12553 4707
rect 12536 4656 12553 4673
rect 12536 4622 12553 4639
rect 12580 4792 12597 4809
rect 12580 4758 12597 4775
rect 12580 4724 12597 4741
rect 12580 4690 12597 4707
rect 12580 4656 12597 4673
rect 12580 4622 12597 4639
rect 12624 4792 12641 4809
rect 12624 4758 12641 4775
rect 12624 4724 12641 4741
rect 12624 4690 12641 4707
rect 12624 4656 12641 4673
rect 12624 4622 12641 4639
rect 13147 4792 13164 4809
rect 13147 4758 13164 4775
rect 13147 4724 13164 4741
rect 13147 4690 13164 4707
rect 13147 4656 13164 4673
rect 13147 4622 13164 4639
rect 13191 4792 13208 4809
rect 13191 4758 13208 4775
rect 13191 4724 13208 4741
rect 13191 4690 13208 4707
rect 13191 4656 13208 4673
rect 13191 4622 13208 4639
rect 13235 4792 13252 4809
rect 13235 4758 13252 4775
rect 13235 4724 13252 4741
rect 13235 4690 13252 4707
rect 13235 4656 13252 4673
rect 13235 4622 13252 4639
rect 13758 4792 13775 4809
rect 13758 4758 13775 4775
rect 13758 4724 13775 4741
rect 13758 4690 13775 4707
rect 13758 4656 13775 4673
rect 13758 4622 13775 4639
rect 13802 4792 13819 4809
rect 13802 4758 13819 4775
rect 13802 4724 13819 4741
rect 13802 4690 13819 4707
rect 13802 4656 13819 4673
rect 13802 4622 13819 4639
rect 13846 4792 13863 4809
rect 13846 4758 13863 4775
rect 13846 4724 13863 4741
rect 13846 4690 13863 4707
rect 13846 4656 13863 4673
rect 13846 4622 13863 4639
rect 14336 4792 14353 4809
rect 14336 4758 14353 4775
rect 14336 4724 14353 4741
rect 14336 4690 14353 4707
rect 14336 4656 14353 4673
rect 14336 4622 14353 4639
rect 14380 4792 14397 4809
rect 14380 4758 14397 4775
rect 14380 4724 14397 4741
rect 14380 4690 14397 4707
rect 14380 4656 14397 4673
rect 14380 4622 14397 4639
rect 14424 4792 14441 4809
rect 14424 4758 14441 4775
rect 14424 4724 14441 4741
rect 14424 4690 14441 4707
rect 14424 4656 14441 4673
rect 14424 4622 14441 4639
rect 14947 4792 14964 4809
rect 14947 4758 14964 4775
rect 14947 4724 14964 4741
rect 14947 4690 14964 4707
rect 14947 4656 14964 4673
rect 14947 4622 14964 4639
rect 14991 4792 15008 4809
rect 14991 4758 15008 4775
rect 14991 4724 15008 4741
rect 14991 4690 15008 4707
rect 14991 4656 15008 4673
rect 14991 4622 15008 4639
rect 15035 4792 15052 4809
rect 15035 4758 15052 4775
rect 15035 4724 15052 4741
rect 15035 4690 15052 4707
rect 15035 4656 15052 4673
rect 15035 4622 15052 4639
rect 15558 4792 15575 4809
rect 15558 4758 15575 4775
rect 15558 4724 15575 4741
rect 15558 4690 15575 4707
rect 15558 4656 15575 4673
rect 15558 4622 15575 4639
rect 15602 4792 15619 4809
rect 15602 4758 15619 4775
rect 15602 4724 15619 4741
rect 15602 4690 15619 4707
rect 15602 4656 15619 4673
rect 15602 4622 15619 4639
rect 15646 4792 15663 4809
rect 15646 4758 15663 4775
rect 15646 4724 15663 4741
rect 15646 4690 15663 4707
rect 15646 4656 15663 4673
rect 15646 4622 15663 4639
<< poly >>
rect 13170 8044 13185 8057
rect 13214 8044 13229 8057
rect 13781 8044 13796 8057
rect 13825 8044 13840 8057
rect 14359 8044 14374 8057
rect 14403 8044 14418 8057
rect 14970 8044 14985 8057
rect 15014 8044 15029 8057
rect 15581 8044 15596 8057
rect 15625 8044 15640 8057
rect 13170 7827 13185 7844
rect 13160 7819 13193 7827
rect 13160 7802 13168 7819
rect 13185 7802 13193 7819
rect 13160 7794 13193 7802
rect 13061 7767 13094 7775
rect 13061 7750 13069 7767
rect 13086 7757 13094 7767
rect 13086 7750 13141 7757
rect 13061 7742 13141 7750
rect 13061 7713 13105 7721
rect 13061 7696 13069 7713
rect 13086 7696 13105 7713
rect 13061 7688 13105 7696
rect 13090 7670 13105 7688
rect 13126 7670 13141 7742
rect 13170 7670 13185 7794
rect 13214 7773 13229 7844
rect 13781 7827 13796 7844
rect 13771 7819 13804 7827
rect 13771 7802 13779 7819
rect 13796 7802 13804 7819
rect 13771 7794 13804 7802
rect 13206 7765 13239 7773
rect 13206 7748 13214 7765
rect 13231 7748 13239 7765
rect 13206 7740 13239 7748
rect 13672 7767 13705 7775
rect 13672 7750 13680 7767
rect 13697 7757 13705 7767
rect 13697 7750 13752 7757
rect 13672 7742 13752 7750
rect 13214 7670 13229 7740
rect 13305 7729 13338 7737
rect 13305 7719 13313 7729
rect 13258 7712 13313 7719
rect 13330 7712 13338 7729
rect 13258 7704 13338 7712
rect 13672 7713 13716 7721
rect 13258 7670 13273 7704
rect 13672 7696 13680 7713
rect 13697 7696 13716 7713
rect 13672 7688 13716 7696
rect 13294 7670 13309 7683
rect 13701 7670 13716 7688
rect 13737 7670 13752 7742
rect 13781 7670 13796 7794
rect 13825 7773 13840 7844
rect 14359 7827 14374 7844
rect 14349 7819 14382 7827
rect 14349 7802 14357 7819
rect 14374 7802 14382 7819
rect 14349 7794 14382 7802
rect 13817 7765 13850 7773
rect 13817 7748 13825 7765
rect 13842 7748 13850 7765
rect 13817 7740 13850 7748
rect 14250 7767 14283 7775
rect 14250 7750 14258 7767
rect 14275 7757 14283 7767
rect 14275 7750 14330 7757
rect 14250 7742 14330 7750
rect 13825 7670 13840 7740
rect 13916 7729 13949 7737
rect 13916 7719 13924 7729
rect 13869 7712 13924 7719
rect 13941 7712 13949 7729
rect 13869 7704 13949 7712
rect 14250 7713 14294 7721
rect 13869 7670 13884 7704
rect 14250 7696 14258 7713
rect 14275 7696 14294 7713
rect 14250 7688 14294 7696
rect 13905 7670 13920 7683
rect 14279 7670 14294 7688
rect 14315 7670 14330 7742
rect 14359 7670 14374 7794
rect 14403 7773 14418 7844
rect 14970 7827 14985 7844
rect 14960 7819 14993 7827
rect 14960 7802 14968 7819
rect 14985 7802 14993 7819
rect 14960 7794 14993 7802
rect 14395 7765 14428 7773
rect 14395 7748 14403 7765
rect 14420 7748 14428 7765
rect 14395 7740 14428 7748
rect 14861 7767 14894 7775
rect 14861 7750 14869 7767
rect 14886 7757 14894 7767
rect 14886 7750 14941 7757
rect 14861 7742 14941 7750
rect 14403 7670 14418 7740
rect 14494 7729 14527 7737
rect 14494 7719 14502 7729
rect 14447 7712 14502 7719
rect 14519 7712 14527 7729
rect 14447 7704 14527 7712
rect 14861 7713 14905 7721
rect 14447 7670 14462 7704
rect 14861 7696 14869 7713
rect 14886 7696 14905 7713
rect 14861 7688 14905 7696
rect 14483 7670 14498 7683
rect 14890 7670 14905 7688
rect 14926 7670 14941 7742
rect 14970 7670 14985 7794
rect 15014 7773 15029 7844
rect 15581 7827 15596 7844
rect 15571 7819 15604 7827
rect 15571 7802 15579 7819
rect 15596 7802 15604 7819
rect 15571 7794 15604 7802
rect 15006 7765 15039 7773
rect 15006 7748 15014 7765
rect 15031 7748 15039 7765
rect 15006 7740 15039 7748
rect 15472 7767 15505 7775
rect 15472 7750 15480 7767
rect 15497 7757 15505 7767
rect 15497 7750 15552 7757
rect 15472 7742 15552 7750
rect 15014 7670 15029 7740
rect 15105 7729 15138 7737
rect 15105 7719 15113 7729
rect 15058 7712 15113 7719
rect 15130 7712 15138 7729
rect 15058 7704 15138 7712
rect 15472 7713 15516 7721
rect 15058 7670 15073 7704
rect 15472 7696 15480 7713
rect 15497 7696 15516 7713
rect 15472 7688 15516 7696
rect 15094 7670 15109 7683
rect 15501 7670 15516 7688
rect 15537 7670 15552 7742
rect 15581 7670 15596 7794
rect 15625 7773 15640 7844
rect 15617 7765 15650 7773
rect 15617 7748 15625 7765
rect 15642 7748 15650 7765
rect 15617 7740 15650 7748
rect 15625 7670 15640 7740
rect 15716 7729 15749 7737
rect 15716 7719 15724 7729
rect 15669 7712 15724 7719
rect 15741 7712 15749 7729
rect 15669 7704 15749 7712
rect 15669 7670 15684 7704
rect 15705 7670 15720 7683
rect 13090 7536 13105 7570
rect 13126 7557 13141 7570
rect 13170 7557 13185 7570
rect 13214 7557 13229 7570
rect 13258 7557 13273 7570
rect 13294 7536 13309 7570
rect 13090 7521 13309 7536
rect 13701 7536 13716 7570
rect 13737 7557 13752 7570
rect 13781 7557 13796 7570
rect 13825 7557 13840 7570
rect 13869 7557 13884 7570
rect 13905 7536 13920 7570
rect 13701 7521 13920 7536
rect 14279 7536 14294 7570
rect 14315 7557 14330 7570
rect 14359 7557 14374 7570
rect 14403 7557 14418 7570
rect 14447 7557 14462 7570
rect 14483 7536 14498 7570
rect 14279 7521 14498 7536
rect 14890 7536 14905 7570
rect 14926 7557 14941 7570
rect 14970 7557 14985 7570
rect 15014 7557 15029 7570
rect 15058 7557 15073 7570
rect 15094 7536 15109 7570
rect 14890 7521 15109 7536
rect 15501 7536 15516 7570
rect 15537 7557 15552 7570
rect 15581 7557 15596 7570
rect 15625 7557 15640 7570
rect 15669 7557 15684 7570
rect 15705 7536 15720 7570
rect 15501 7521 15720 7536
rect 12559 7394 12574 7407
rect 12603 7394 12618 7407
rect 13170 7394 13185 7407
rect 13214 7394 13229 7407
rect 13781 7394 13796 7407
rect 13825 7394 13840 7407
rect 14359 7394 14374 7407
rect 14403 7394 14418 7407
rect 14970 7394 14985 7407
rect 15014 7394 15029 7407
rect 15581 7394 15596 7407
rect 15625 7394 15640 7407
rect 12559 7177 12574 7194
rect 12549 7169 12582 7177
rect 12549 7152 12557 7169
rect 12574 7152 12582 7169
rect 12549 7144 12582 7152
rect 12450 7117 12483 7125
rect 12450 7100 12458 7117
rect 12475 7107 12483 7117
rect 12475 7100 12530 7107
rect 12450 7092 12530 7100
rect 12450 7063 12494 7071
rect 12450 7046 12458 7063
rect 12475 7046 12494 7063
rect 12450 7038 12494 7046
rect 12479 7020 12494 7038
rect 12515 7020 12530 7092
rect 12559 7020 12574 7144
rect 12603 7123 12618 7194
rect 13170 7177 13185 7194
rect 13160 7169 13193 7177
rect 13160 7152 13168 7169
rect 13185 7152 13193 7169
rect 13160 7144 13193 7152
rect 12595 7115 12628 7123
rect 12595 7098 12603 7115
rect 12620 7098 12628 7115
rect 12595 7090 12628 7098
rect 13061 7117 13094 7125
rect 13061 7100 13069 7117
rect 13086 7107 13094 7117
rect 13086 7100 13141 7107
rect 13061 7092 13141 7100
rect 12603 7020 12618 7090
rect 12694 7079 12727 7087
rect 12694 7069 12702 7079
rect 12647 7062 12702 7069
rect 12719 7062 12727 7079
rect 12647 7054 12727 7062
rect 13061 7063 13105 7071
rect 12647 7020 12662 7054
rect 13061 7046 13069 7063
rect 13086 7046 13105 7063
rect 13061 7038 13105 7046
rect 12683 7020 12698 7033
rect 13090 7020 13105 7038
rect 13126 7020 13141 7092
rect 13170 7020 13185 7144
rect 13214 7123 13229 7194
rect 13781 7177 13796 7194
rect 13771 7169 13804 7177
rect 13771 7152 13779 7169
rect 13796 7152 13804 7169
rect 13771 7144 13804 7152
rect 13206 7115 13239 7123
rect 13206 7098 13214 7115
rect 13231 7098 13239 7115
rect 13206 7090 13239 7098
rect 13672 7117 13705 7125
rect 13672 7100 13680 7117
rect 13697 7107 13705 7117
rect 13697 7100 13752 7107
rect 13672 7092 13752 7100
rect 13214 7020 13229 7090
rect 13305 7079 13338 7087
rect 13305 7069 13313 7079
rect 13258 7062 13313 7069
rect 13330 7062 13338 7079
rect 13258 7054 13338 7062
rect 13672 7063 13716 7071
rect 13258 7020 13273 7054
rect 13672 7046 13680 7063
rect 13697 7046 13716 7063
rect 13672 7038 13716 7046
rect 13294 7020 13309 7033
rect 13701 7020 13716 7038
rect 13737 7020 13752 7092
rect 13781 7020 13796 7144
rect 13825 7123 13840 7194
rect 14359 7177 14374 7194
rect 14349 7169 14382 7177
rect 14349 7152 14357 7169
rect 14374 7152 14382 7169
rect 14349 7144 14382 7152
rect 13817 7115 13850 7123
rect 13817 7098 13825 7115
rect 13842 7098 13850 7115
rect 13817 7090 13850 7098
rect 14250 7117 14283 7125
rect 14250 7100 14258 7117
rect 14275 7107 14283 7117
rect 14275 7100 14330 7107
rect 14250 7092 14330 7100
rect 13825 7020 13840 7090
rect 13916 7079 13949 7087
rect 13916 7069 13924 7079
rect 13869 7062 13924 7069
rect 13941 7062 13949 7079
rect 13869 7054 13949 7062
rect 14250 7063 14294 7071
rect 13869 7020 13884 7054
rect 14250 7046 14258 7063
rect 14275 7046 14294 7063
rect 14250 7038 14294 7046
rect 13905 7020 13920 7033
rect 14279 7020 14294 7038
rect 14315 7020 14330 7092
rect 14359 7020 14374 7144
rect 14403 7123 14418 7194
rect 14970 7177 14985 7194
rect 14960 7169 14993 7177
rect 14960 7152 14968 7169
rect 14985 7152 14993 7169
rect 14960 7144 14993 7152
rect 14395 7115 14428 7123
rect 14395 7098 14403 7115
rect 14420 7098 14428 7115
rect 14395 7090 14428 7098
rect 14861 7117 14894 7125
rect 14861 7100 14869 7117
rect 14886 7107 14894 7117
rect 14886 7100 14941 7107
rect 14861 7092 14941 7100
rect 14403 7020 14418 7090
rect 14494 7079 14527 7087
rect 14494 7069 14502 7079
rect 14447 7062 14502 7069
rect 14519 7062 14527 7079
rect 14447 7054 14527 7062
rect 14861 7063 14905 7071
rect 14447 7020 14462 7054
rect 14861 7046 14869 7063
rect 14886 7046 14905 7063
rect 14861 7038 14905 7046
rect 14483 7020 14498 7033
rect 14890 7020 14905 7038
rect 14926 7020 14941 7092
rect 14970 7020 14985 7144
rect 15014 7123 15029 7194
rect 15581 7177 15596 7194
rect 15571 7169 15604 7177
rect 15571 7152 15579 7169
rect 15596 7152 15604 7169
rect 15571 7144 15604 7152
rect 15006 7115 15039 7123
rect 15006 7098 15014 7115
rect 15031 7098 15039 7115
rect 15006 7090 15039 7098
rect 15472 7117 15505 7125
rect 15472 7100 15480 7117
rect 15497 7107 15505 7117
rect 15497 7100 15552 7107
rect 15472 7092 15552 7100
rect 15014 7020 15029 7090
rect 15105 7079 15138 7087
rect 15105 7069 15113 7079
rect 15058 7062 15113 7069
rect 15130 7062 15138 7079
rect 15058 7054 15138 7062
rect 15472 7063 15516 7071
rect 15058 7020 15073 7054
rect 15472 7046 15480 7063
rect 15497 7046 15516 7063
rect 15472 7038 15516 7046
rect 15094 7020 15109 7033
rect 15501 7020 15516 7038
rect 15537 7020 15552 7092
rect 15581 7020 15596 7144
rect 15625 7123 15640 7194
rect 15617 7115 15650 7123
rect 15617 7098 15625 7115
rect 15642 7098 15650 7115
rect 15617 7090 15650 7098
rect 15625 7020 15640 7090
rect 15716 7079 15749 7087
rect 15716 7069 15724 7079
rect 15669 7062 15724 7069
rect 15741 7062 15749 7079
rect 15669 7054 15749 7062
rect 15669 7020 15684 7054
rect 15705 7020 15720 7033
rect 12479 6886 12494 6920
rect 12515 6907 12530 6920
rect 12559 6907 12574 6920
rect 12603 6907 12618 6920
rect 12647 6907 12662 6920
rect 12683 6886 12698 6920
rect 12479 6871 12698 6886
rect 13090 6886 13105 6920
rect 13126 6907 13141 6920
rect 13170 6907 13185 6920
rect 13214 6907 13229 6920
rect 13258 6907 13273 6920
rect 13294 6886 13309 6920
rect 13090 6871 13309 6886
rect 13701 6886 13716 6920
rect 13737 6907 13752 6920
rect 13781 6907 13796 6920
rect 13825 6907 13840 6920
rect 13869 6907 13884 6920
rect 13905 6886 13920 6920
rect 13701 6871 13920 6886
rect 14279 6886 14294 6920
rect 14315 6907 14330 6920
rect 14359 6907 14374 6920
rect 14403 6907 14418 6920
rect 14447 6907 14462 6920
rect 14483 6886 14498 6920
rect 14279 6871 14498 6886
rect 14890 6886 14905 6920
rect 14926 6907 14941 6920
rect 14970 6907 14985 6920
rect 15014 6907 15029 6920
rect 15058 6907 15073 6920
rect 15094 6886 15109 6920
rect 14890 6871 15109 6886
rect 15501 6886 15516 6920
rect 15537 6907 15552 6920
rect 15581 6907 15596 6920
rect 15625 6907 15640 6920
rect 15669 6907 15684 6920
rect 15705 6886 15720 6920
rect 15501 6871 15720 6886
rect 12559 6754 12574 6767
rect 12603 6754 12618 6767
rect 13170 6754 13185 6767
rect 13214 6754 13229 6767
rect 13781 6754 13796 6767
rect 13825 6754 13840 6767
rect 14359 6754 14374 6767
rect 14403 6754 14418 6767
rect 14970 6754 14985 6767
rect 15014 6754 15029 6767
rect 15581 6754 15596 6767
rect 15625 6754 15640 6767
rect 12559 6537 12574 6554
rect 12549 6529 12582 6537
rect 12549 6512 12557 6529
rect 12574 6512 12582 6529
rect 12549 6504 12582 6512
rect 12450 6477 12483 6485
rect 12450 6460 12458 6477
rect 12475 6467 12483 6477
rect 12475 6460 12530 6467
rect 12450 6452 12530 6460
rect 12450 6423 12494 6431
rect 12450 6406 12458 6423
rect 12475 6406 12494 6423
rect 12450 6398 12494 6406
rect 12479 6380 12494 6398
rect 12515 6380 12530 6452
rect 12559 6380 12574 6504
rect 12603 6483 12618 6554
rect 13170 6537 13185 6554
rect 13160 6529 13193 6537
rect 13160 6512 13168 6529
rect 13185 6512 13193 6529
rect 13160 6504 13193 6512
rect 12595 6475 12628 6483
rect 12595 6458 12603 6475
rect 12620 6458 12628 6475
rect 12595 6450 12628 6458
rect 13061 6477 13094 6485
rect 13061 6460 13069 6477
rect 13086 6467 13094 6477
rect 13086 6460 13141 6467
rect 13061 6452 13141 6460
rect 12603 6380 12618 6450
rect 12694 6439 12727 6447
rect 12694 6429 12702 6439
rect 12647 6422 12702 6429
rect 12719 6422 12727 6439
rect 12647 6414 12727 6422
rect 13061 6423 13105 6431
rect 12647 6380 12662 6414
rect 13061 6406 13069 6423
rect 13086 6406 13105 6423
rect 13061 6398 13105 6406
rect 12683 6380 12698 6393
rect 13090 6380 13105 6398
rect 13126 6380 13141 6452
rect 13170 6380 13185 6504
rect 13214 6483 13229 6554
rect 13781 6537 13796 6554
rect 13771 6529 13804 6537
rect 13771 6512 13779 6529
rect 13796 6512 13804 6529
rect 13771 6504 13804 6512
rect 13206 6475 13239 6483
rect 13206 6458 13214 6475
rect 13231 6458 13239 6475
rect 13206 6450 13239 6458
rect 13672 6477 13705 6485
rect 13672 6460 13680 6477
rect 13697 6467 13705 6477
rect 13697 6460 13752 6467
rect 13672 6452 13752 6460
rect 13214 6380 13229 6450
rect 13305 6439 13338 6447
rect 13305 6429 13313 6439
rect 13258 6422 13313 6429
rect 13330 6422 13338 6439
rect 13258 6414 13338 6422
rect 13672 6423 13716 6431
rect 13258 6380 13273 6414
rect 13672 6406 13680 6423
rect 13697 6406 13716 6423
rect 13672 6398 13716 6406
rect 13294 6380 13309 6393
rect 13701 6380 13716 6398
rect 13737 6380 13752 6452
rect 13781 6380 13796 6504
rect 13825 6483 13840 6554
rect 14359 6537 14374 6554
rect 14349 6529 14382 6537
rect 14349 6512 14357 6529
rect 14374 6512 14382 6529
rect 14349 6504 14382 6512
rect 13817 6475 13850 6483
rect 13817 6458 13825 6475
rect 13842 6458 13850 6475
rect 13817 6450 13850 6458
rect 14250 6477 14283 6485
rect 14250 6460 14258 6477
rect 14275 6467 14283 6477
rect 14275 6460 14330 6467
rect 14250 6452 14330 6460
rect 13825 6380 13840 6450
rect 13916 6439 13949 6447
rect 13916 6429 13924 6439
rect 13869 6422 13924 6429
rect 13941 6422 13949 6439
rect 13869 6414 13949 6422
rect 14250 6423 14294 6431
rect 13869 6380 13884 6414
rect 14250 6406 14258 6423
rect 14275 6406 14294 6423
rect 14250 6398 14294 6406
rect 13905 6380 13920 6393
rect 14279 6380 14294 6398
rect 14315 6380 14330 6452
rect 14359 6380 14374 6504
rect 14403 6483 14418 6554
rect 14970 6537 14985 6554
rect 14960 6529 14993 6537
rect 14960 6512 14968 6529
rect 14985 6512 14993 6529
rect 14960 6504 14993 6512
rect 14395 6475 14428 6483
rect 14395 6458 14403 6475
rect 14420 6458 14428 6475
rect 14395 6450 14428 6458
rect 14861 6477 14894 6485
rect 14861 6460 14869 6477
rect 14886 6467 14894 6477
rect 14886 6460 14941 6467
rect 14861 6452 14941 6460
rect 14403 6380 14418 6450
rect 14494 6439 14527 6447
rect 14494 6429 14502 6439
rect 14447 6422 14502 6429
rect 14519 6422 14527 6439
rect 14447 6414 14527 6422
rect 14861 6423 14905 6431
rect 14447 6380 14462 6414
rect 14861 6406 14869 6423
rect 14886 6406 14905 6423
rect 14861 6398 14905 6406
rect 14483 6380 14498 6393
rect 14890 6380 14905 6398
rect 14926 6380 14941 6452
rect 14970 6380 14985 6504
rect 15014 6483 15029 6554
rect 15581 6537 15596 6554
rect 15571 6529 15604 6537
rect 15571 6512 15579 6529
rect 15596 6512 15604 6529
rect 15571 6504 15604 6512
rect 15006 6475 15039 6483
rect 15006 6458 15014 6475
rect 15031 6458 15039 6475
rect 15006 6450 15039 6458
rect 15472 6477 15505 6485
rect 15472 6460 15480 6477
rect 15497 6467 15505 6477
rect 15497 6460 15552 6467
rect 15472 6452 15552 6460
rect 15014 6380 15029 6450
rect 15105 6439 15138 6447
rect 15105 6429 15113 6439
rect 15058 6422 15113 6429
rect 15130 6422 15138 6439
rect 15058 6414 15138 6422
rect 15472 6423 15516 6431
rect 15058 6380 15073 6414
rect 15472 6406 15480 6423
rect 15497 6406 15516 6423
rect 15472 6398 15516 6406
rect 15094 6380 15109 6393
rect 15501 6380 15516 6398
rect 15537 6380 15552 6452
rect 15581 6380 15596 6504
rect 15625 6483 15640 6554
rect 15617 6475 15650 6483
rect 15617 6458 15625 6475
rect 15642 6458 15650 6475
rect 15617 6450 15650 6458
rect 15625 6380 15640 6450
rect 15716 6439 15749 6447
rect 15716 6429 15724 6439
rect 15669 6422 15724 6429
rect 15741 6422 15749 6439
rect 15669 6414 15749 6422
rect 15669 6380 15684 6414
rect 15705 6380 15720 6393
rect 12479 6246 12494 6280
rect 12515 6267 12530 6280
rect 12559 6267 12574 6280
rect 12603 6267 12618 6280
rect 12647 6267 12662 6280
rect 12683 6246 12698 6280
rect 12479 6231 12698 6246
rect 13090 6246 13105 6280
rect 13126 6267 13141 6280
rect 13170 6267 13185 6280
rect 13214 6267 13229 6280
rect 13258 6267 13273 6280
rect 13294 6246 13309 6280
rect 13090 6231 13309 6246
rect 13701 6246 13716 6280
rect 13737 6267 13752 6280
rect 13781 6267 13796 6280
rect 13825 6267 13840 6280
rect 13869 6267 13884 6280
rect 13905 6246 13920 6280
rect 13701 6231 13920 6246
rect 14279 6246 14294 6280
rect 14315 6267 14330 6280
rect 14359 6267 14374 6280
rect 14403 6267 14418 6280
rect 14447 6267 14462 6280
rect 14483 6246 14498 6280
rect 14279 6231 14498 6246
rect 14890 6246 14905 6280
rect 14926 6267 14941 6280
rect 14970 6267 14985 6280
rect 15014 6267 15029 6280
rect 15058 6267 15073 6280
rect 15094 6246 15109 6280
rect 14890 6231 15109 6246
rect 15501 6246 15516 6280
rect 15537 6267 15552 6280
rect 15581 6267 15596 6280
rect 15625 6267 15640 6280
rect 15669 6267 15684 6280
rect 15705 6246 15720 6280
rect 15501 6231 15720 6246
rect 12559 6104 12574 6117
rect 12603 6104 12618 6117
rect 13170 6104 13185 6117
rect 13214 6104 13229 6117
rect 13781 6104 13796 6117
rect 13825 6104 13840 6117
rect 14359 6104 14374 6117
rect 14403 6104 14418 6117
rect 14970 6104 14985 6117
rect 15014 6104 15029 6117
rect 15581 6104 15596 6117
rect 15625 6104 15640 6117
rect 12559 5887 12574 5904
rect 12549 5879 12582 5887
rect 12549 5862 12557 5879
rect 12574 5862 12582 5879
rect 12549 5854 12582 5862
rect 12450 5827 12483 5835
rect 12450 5810 12458 5827
rect 12475 5817 12483 5827
rect 12475 5810 12530 5817
rect 12450 5802 12530 5810
rect 12450 5773 12494 5781
rect 12450 5756 12458 5773
rect 12475 5756 12494 5773
rect 12450 5748 12494 5756
rect 12479 5730 12494 5748
rect 12515 5730 12530 5802
rect 12559 5730 12574 5854
rect 12603 5833 12618 5904
rect 13170 5887 13185 5904
rect 13160 5879 13193 5887
rect 13160 5862 13168 5879
rect 13185 5862 13193 5879
rect 13160 5854 13193 5862
rect 12595 5825 12628 5833
rect 12595 5808 12603 5825
rect 12620 5808 12628 5825
rect 12595 5800 12628 5808
rect 13061 5827 13094 5835
rect 13061 5810 13069 5827
rect 13086 5817 13094 5827
rect 13086 5810 13141 5817
rect 13061 5802 13141 5810
rect 12603 5730 12618 5800
rect 12694 5789 12727 5797
rect 12694 5779 12702 5789
rect 12647 5772 12702 5779
rect 12719 5772 12727 5789
rect 12647 5764 12727 5772
rect 13061 5773 13105 5781
rect 12647 5730 12662 5764
rect 13061 5756 13069 5773
rect 13086 5756 13105 5773
rect 13061 5748 13105 5756
rect 12683 5730 12698 5743
rect 13090 5730 13105 5748
rect 13126 5730 13141 5802
rect 13170 5730 13185 5854
rect 13214 5833 13229 5904
rect 13781 5887 13796 5904
rect 13771 5879 13804 5887
rect 13771 5862 13779 5879
rect 13796 5862 13804 5879
rect 13771 5854 13804 5862
rect 13206 5825 13239 5833
rect 13206 5808 13214 5825
rect 13231 5808 13239 5825
rect 13206 5800 13239 5808
rect 13672 5827 13705 5835
rect 13672 5810 13680 5827
rect 13697 5817 13705 5827
rect 13697 5810 13752 5817
rect 13672 5802 13752 5810
rect 13214 5730 13229 5800
rect 13305 5789 13338 5797
rect 13305 5779 13313 5789
rect 13258 5772 13313 5779
rect 13330 5772 13338 5789
rect 13258 5764 13338 5772
rect 13672 5773 13716 5781
rect 13258 5730 13273 5764
rect 13672 5756 13680 5773
rect 13697 5756 13716 5773
rect 13672 5748 13716 5756
rect 13294 5730 13309 5743
rect 13701 5730 13716 5748
rect 13737 5730 13752 5802
rect 13781 5730 13796 5854
rect 13825 5833 13840 5904
rect 14359 5887 14374 5904
rect 14349 5879 14382 5887
rect 14349 5862 14357 5879
rect 14374 5862 14382 5879
rect 14349 5854 14382 5862
rect 13817 5825 13850 5833
rect 13817 5808 13825 5825
rect 13842 5808 13850 5825
rect 13817 5800 13850 5808
rect 14250 5827 14283 5835
rect 14250 5810 14258 5827
rect 14275 5817 14283 5827
rect 14275 5810 14330 5817
rect 14250 5802 14330 5810
rect 13825 5730 13840 5800
rect 13916 5789 13949 5797
rect 13916 5779 13924 5789
rect 13869 5772 13924 5779
rect 13941 5772 13949 5789
rect 13869 5764 13949 5772
rect 14250 5773 14294 5781
rect 13869 5730 13884 5764
rect 14250 5756 14258 5773
rect 14275 5756 14294 5773
rect 14250 5748 14294 5756
rect 13905 5730 13920 5743
rect 14279 5730 14294 5748
rect 14315 5730 14330 5802
rect 14359 5730 14374 5854
rect 14403 5833 14418 5904
rect 14970 5887 14985 5904
rect 14960 5879 14993 5887
rect 14960 5862 14968 5879
rect 14985 5862 14993 5879
rect 14960 5854 14993 5862
rect 14395 5825 14428 5833
rect 14395 5808 14403 5825
rect 14420 5808 14428 5825
rect 14395 5800 14428 5808
rect 14861 5827 14894 5835
rect 14861 5810 14869 5827
rect 14886 5817 14894 5827
rect 14886 5810 14941 5817
rect 14861 5802 14941 5810
rect 14403 5730 14418 5800
rect 14494 5789 14527 5797
rect 14494 5779 14502 5789
rect 14447 5772 14502 5779
rect 14519 5772 14527 5789
rect 14447 5764 14527 5772
rect 14861 5773 14905 5781
rect 14447 5730 14462 5764
rect 14861 5756 14869 5773
rect 14886 5756 14905 5773
rect 14861 5748 14905 5756
rect 14483 5730 14498 5743
rect 14890 5730 14905 5748
rect 14926 5730 14941 5802
rect 14970 5730 14985 5854
rect 15014 5833 15029 5904
rect 15581 5887 15596 5904
rect 15571 5879 15604 5887
rect 15571 5862 15579 5879
rect 15596 5862 15604 5879
rect 15571 5854 15604 5862
rect 15006 5825 15039 5833
rect 15006 5808 15014 5825
rect 15031 5808 15039 5825
rect 15006 5800 15039 5808
rect 15472 5827 15505 5835
rect 15472 5810 15480 5827
rect 15497 5817 15505 5827
rect 15497 5810 15552 5817
rect 15472 5802 15552 5810
rect 15014 5730 15029 5800
rect 15105 5789 15138 5797
rect 15105 5779 15113 5789
rect 15058 5772 15113 5779
rect 15130 5772 15138 5789
rect 15058 5764 15138 5772
rect 15472 5773 15516 5781
rect 15058 5730 15073 5764
rect 15472 5756 15480 5773
rect 15497 5756 15516 5773
rect 15472 5748 15516 5756
rect 15094 5730 15109 5743
rect 15501 5730 15516 5748
rect 15537 5730 15552 5802
rect 15581 5730 15596 5854
rect 15625 5833 15640 5904
rect 15617 5825 15650 5833
rect 15617 5808 15625 5825
rect 15642 5808 15650 5825
rect 15617 5800 15650 5808
rect 15625 5730 15640 5800
rect 15716 5789 15749 5797
rect 15716 5779 15724 5789
rect 15669 5772 15724 5779
rect 15741 5772 15749 5789
rect 15669 5764 15749 5772
rect 15669 5730 15684 5764
rect 15705 5730 15720 5743
rect 12479 5596 12494 5630
rect 12515 5617 12530 5630
rect 12559 5617 12574 5630
rect 12603 5617 12618 5630
rect 12647 5617 12662 5630
rect 12683 5596 12698 5630
rect 12479 5581 12698 5596
rect 13090 5596 13105 5630
rect 13126 5617 13141 5630
rect 13170 5617 13185 5630
rect 13214 5617 13229 5630
rect 13258 5617 13273 5630
rect 13294 5596 13309 5630
rect 13090 5581 13309 5596
rect 13701 5596 13716 5630
rect 13737 5617 13752 5630
rect 13781 5617 13796 5630
rect 13825 5617 13840 5630
rect 13869 5617 13884 5630
rect 13905 5596 13920 5630
rect 13701 5581 13920 5596
rect 14279 5596 14294 5630
rect 14315 5617 14330 5630
rect 14359 5617 14374 5630
rect 14403 5617 14418 5630
rect 14447 5617 14462 5630
rect 14483 5596 14498 5630
rect 14279 5581 14498 5596
rect 14890 5596 14905 5630
rect 14926 5617 14941 5630
rect 14970 5617 14985 5630
rect 15014 5617 15029 5630
rect 15058 5617 15073 5630
rect 15094 5596 15109 5630
rect 14890 5581 15109 5596
rect 15501 5596 15516 5630
rect 15537 5617 15552 5630
rect 15581 5617 15596 5630
rect 15625 5617 15640 5630
rect 15669 5617 15684 5630
rect 15705 5596 15720 5630
rect 15501 5581 15720 5596
rect 12559 5454 12574 5467
rect 12603 5454 12618 5467
rect 13170 5454 13185 5467
rect 13214 5454 13229 5467
rect 13781 5454 13796 5467
rect 13825 5454 13840 5467
rect 14359 5454 14374 5467
rect 14403 5454 14418 5467
rect 14970 5454 14985 5467
rect 15014 5454 15029 5467
rect 15581 5454 15596 5467
rect 15625 5454 15640 5467
rect 12559 5237 12574 5254
rect 12549 5229 12582 5237
rect 12549 5212 12557 5229
rect 12574 5212 12582 5229
rect 12549 5204 12582 5212
rect 12450 5177 12483 5185
rect 12450 5160 12458 5177
rect 12475 5167 12483 5177
rect 12475 5160 12530 5167
rect 12450 5152 12530 5160
rect 12450 5123 12494 5131
rect 12450 5106 12458 5123
rect 12475 5106 12494 5123
rect 12450 5098 12494 5106
rect 12479 5080 12494 5098
rect 12515 5080 12530 5152
rect 12559 5080 12574 5204
rect 12603 5183 12618 5254
rect 13170 5237 13185 5254
rect 13160 5229 13193 5237
rect 13160 5212 13168 5229
rect 13185 5212 13193 5229
rect 13160 5204 13193 5212
rect 12595 5175 12628 5183
rect 12595 5158 12603 5175
rect 12620 5158 12628 5175
rect 12595 5150 12628 5158
rect 13061 5177 13094 5185
rect 13061 5160 13069 5177
rect 13086 5167 13094 5177
rect 13086 5160 13141 5167
rect 13061 5152 13141 5160
rect 12603 5080 12618 5150
rect 12694 5139 12727 5147
rect 12694 5129 12702 5139
rect 12647 5122 12702 5129
rect 12719 5122 12727 5139
rect 12647 5114 12727 5122
rect 13061 5123 13105 5131
rect 12647 5080 12662 5114
rect 13061 5106 13069 5123
rect 13086 5106 13105 5123
rect 13061 5098 13105 5106
rect 12683 5080 12698 5093
rect 13090 5080 13105 5098
rect 13126 5080 13141 5152
rect 13170 5080 13185 5204
rect 13214 5183 13229 5254
rect 13781 5237 13796 5254
rect 13771 5229 13804 5237
rect 13771 5212 13779 5229
rect 13796 5212 13804 5229
rect 13771 5204 13804 5212
rect 13206 5175 13239 5183
rect 13206 5158 13214 5175
rect 13231 5158 13239 5175
rect 13206 5150 13239 5158
rect 13672 5177 13705 5185
rect 13672 5160 13680 5177
rect 13697 5167 13705 5177
rect 13697 5160 13752 5167
rect 13672 5152 13752 5160
rect 13214 5080 13229 5150
rect 13305 5139 13338 5147
rect 13305 5129 13313 5139
rect 13258 5122 13313 5129
rect 13330 5122 13338 5139
rect 13258 5114 13338 5122
rect 13672 5123 13716 5131
rect 13258 5080 13273 5114
rect 13672 5106 13680 5123
rect 13697 5106 13716 5123
rect 13672 5098 13716 5106
rect 13294 5080 13309 5093
rect 13701 5080 13716 5098
rect 13737 5080 13752 5152
rect 13781 5080 13796 5204
rect 13825 5183 13840 5254
rect 14359 5237 14374 5254
rect 14349 5229 14382 5237
rect 14349 5212 14357 5229
rect 14374 5212 14382 5229
rect 14349 5204 14382 5212
rect 13817 5175 13850 5183
rect 13817 5158 13825 5175
rect 13842 5158 13850 5175
rect 13817 5150 13850 5158
rect 14250 5177 14283 5185
rect 14250 5160 14258 5177
rect 14275 5167 14283 5177
rect 14275 5160 14330 5167
rect 14250 5152 14330 5160
rect 13825 5080 13840 5150
rect 13916 5139 13949 5147
rect 13916 5129 13924 5139
rect 13869 5122 13924 5129
rect 13941 5122 13949 5139
rect 13869 5114 13949 5122
rect 14250 5123 14294 5131
rect 13869 5080 13884 5114
rect 14250 5106 14258 5123
rect 14275 5106 14294 5123
rect 14250 5098 14294 5106
rect 13905 5080 13920 5093
rect 14279 5080 14294 5098
rect 14315 5080 14330 5152
rect 14359 5080 14374 5204
rect 14403 5183 14418 5254
rect 14970 5237 14985 5254
rect 14960 5229 14993 5237
rect 14960 5212 14968 5229
rect 14985 5212 14993 5229
rect 14960 5204 14993 5212
rect 14395 5175 14428 5183
rect 14395 5158 14403 5175
rect 14420 5158 14428 5175
rect 14395 5150 14428 5158
rect 14861 5177 14894 5185
rect 14861 5160 14869 5177
rect 14886 5167 14894 5177
rect 14886 5160 14941 5167
rect 14861 5152 14941 5160
rect 14403 5080 14418 5150
rect 14494 5139 14527 5147
rect 14494 5129 14502 5139
rect 14447 5122 14502 5129
rect 14519 5122 14527 5139
rect 14447 5114 14527 5122
rect 14861 5123 14905 5131
rect 14447 5080 14462 5114
rect 14861 5106 14869 5123
rect 14886 5106 14905 5123
rect 14861 5098 14905 5106
rect 14483 5080 14498 5093
rect 14890 5080 14905 5098
rect 14926 5080 14941 5152
rect 14970 5080 14985 5204
rect 15014 5183 15029 5254
rect 15581 5237 15596 5254
rect 15571 5229 15604 5237
rect 15571 5212 15579 5229
rect 15596 5212 15604 5229
rect 15571 5204 15604 5212
rect 15006 5175 15039 5183
rect 15006 5158 15014 5175
rect 15031 5158 15039 5175
rect 15006 5150 15039 5158
rect 15472 5177 15505 5185
rect 15472 5160 15480 5177
rect 15497 5167 15505 5177
rect 15497 5160 15552 5167
rect 15472 5152 15552 5160
rect 15014 5080 15029 5150
rect 15105 5139 15138 5147
rect 15105 5129 15113 5139
rect 15058 5122 15113 5129
rect 15130 5122 15138 5139
rect 15058 5114 15138 5122
rect 15472 5123 15516 5131
rect 15058 5080 15073 5114
rect 15472 5106 15480 5123
rect 15497 5106 15516 5123
rect 15472 5098 15516 5106
rect 15094 5080 15109 5093
rect 15501 5080 15516 5098
rect 15537 5080 15552 5152
rect 15581 5080 15596 5204
rect 15625 5183 15640 5254
rect 15617 5175 15650 5183
rect 15617 5158 15625 5175
rect 15642 5158 15650 5175
rect 15617 5150 15650 5158
rect 15625 5080 15640 5150
rect 15716 5139 15749 5147
rect 15716 5129 15724 5139
rect 15669 5122 15724 5129
rect 15741 5122 15749 5139
rect 15669 5114 15749 5122
rect 15669 5080 15684 5114
rect 15705 5080 15720 5093
rect 12479 4946 12494 4980
rect 12515 4967 12530 4980
rect 12559 4967 12574 4980
rect 12603 4967 12618 4980
rect 12647 4967 12662 4980
rect 12683 4946 12698 4980
rect 12479 4931 12698 4946
rect 13090 4946 13105 4980
rect 13126 4967 13141 4980
rect 13170 4967 13185 4980
rect 13214 4967 13229 4980
rect 13258 4967 13273 4980
rect 13294 4946 13309 4980
rect 13090 4931 13309 4946
rect 13701 4946 13716 4980
rect 13737 4967 13752 4980
rect 13781 4967 13796 4980
rect 13825 4967 13840 4980
rect 13869 4967 13884 4980
rect 13905 4946 13920 4980
rect 13701 4931 13920 4946
rect 14279 4946 14294 4980
rect 14315 4967 14330 4980
rect 14359 4967 14374 4980
rect 14403 4967 14418 4980
rect 14447 4967 14462 4980
rect 14483 4946 14498 4980
rect 14279 4931 14498 4946
rect 14890 4946 14905 4980
rect 14926 4967 14941 4980
rect 14970 4967 14985 4980
rect 15014 4967 15029 4980
rect 15058 4967 15073 4980
rect 15094 4946 15109 4980
rect 14890 4931 15109 4946
rect 15501 4946 15516 4980
rect 15537 4967 15552 4980
rect 15581 4967 15596 4980
rect 15625 4967 15640 4980
rect 15669 4967 15684 4980
rect 15705 4946 15720 4980
rect 15501 4931 15720 4946
rect 12559 4814 12574 4827
rect 12603 4814 12618 4827
rect 13170 4814 13185 4827
rect 13214 4814 13229 4827
rect 13781 4814 13796 4827
rect 13825 4814 13840 4827
rect 14359 4814 14374 4827
rect 14403 4814 14418 4827
rect 14970 4814 14985 4827
rect 15014 4814 15029 4827
rect 15581 4814 15596 4827
rect 15625 4814 15640 4827
rect 12559 4597 12574 4614
rect 12549 4589 12582 4597
rect 12549 4572 12557 4589
rect 12574 4572 12582 4589
rect 12549 4564 12582 4572
rect 12450 4537 12483 4545
rect 12450 4520 12458 4537
rect 12475 4527 12483 4537
rect 12475 4520 12530 4527
rect 12450 4512 12530 4520
rect 12450 4483 12494 4491
rect 12450 4466 12458 4483
rect 12475 4466 12494 4483
rect 12450 4458 12494 4466
rect 12479 4440 12494 4458
rect 12515 4440 12530 4512
rect 12559 4440 12574 4564
rect 12603 4543 12618 4614
rect 13170 4597 13185 4614
rect 13160 4589 13193 4597
rect 13160 4572 13168 4589
rect 13185 4572 13193 4589
rect 13160 4564 13193 4572
rect 12595 4535 12628 4543
rect 12595 4518 12603 4535
rect 12620 4518 12628 4535
rect 12595 4510 12628 4518
rect 13061 4537 13094 4545
rect 13061 4520 13069 4537
rect 13086 4527 13094 4537
rect 13086 4520 13141 4527
rect 13061 4512 13141 4520
rect 12603 4440 12618 4510
rect 12694 4499 12727 4507
rect 12694 4489 12702 4499
rect 12647 4482 12702 4489
rect 12719 4482 12727 4499
rect 12647 4474 12727 4482
rect 13061 4483 13105 4491
rect 12647 4440 12662 4474
rect 13061 4466 13069 4483
rect 13086 4466 13105 4483
rect 13061 4458 13105 4466
rect 12683 4440 12698 4453
rect 13090 4440 13105 4458
rect 13126 4440 13141 4512
rect 13170 4440 13185 4564
rect 13214 4543 13229 4614
rect 13781 4597 13796 4614
rect 13771 4589 13804 4597
rect 13771 4572 13779 4589
rect 13796 4572 13804 4589
rect 13771 4564 13804 4572
rect 13206 4535 13239 4543
rect 13206 4518 13214 4535
rect 13231 4518 13239 4535
rect 13206 4510 13239 4518
rect 13672 4537 13705 4545
rect 13672 4520 13680 4537
rect 13697 4527 13705 4537
rect 13697 4520 13752 4527
rect 13672 4512 13752 4520
rect 13214 4440 13229 4510
rect 13305 4499 13338 4507
rect 13305 4489 13313 4499
rect 13258 4482 13313 4489
rect 13330 4482 13338 4499
rect 13258 4474 13338 4482
rect 13672 4483 13716 4491
rect 13258 4440 13273 4474
rect 13672 4466 13680 4483
rect 13697 4466 13716 4483
rect 13672 4458 13716 4466
rect 13294 4440 13309 4453
rect 13701 4440 13716 4458
rect 13737 4440 13752 4512
rect 13781 4440 13796 4564
rect 13825 4543 13840 4614
rect 14359 4597 14374 4614
rect 14349 4589 14382 4597
rect 14349 4572 14357 4589
rect 14374 4572 14382 4589
rect 14349 4564 14382 4572
rect 13817 4535 13850 4543
rect 13817 4518 13825 4535
rect 13842 4518 13850 4535
rect 13817 4510 13850 4518
rect 14250 4537 14283 4545
rect 14250 4520 14258 4537
rect 14275 4527 14283 4537
rect 14275 4520 14330 4527
rect 14250 4512 14330 4520
rect 13825 4440 13840 4510
rect 13916 4499 13949 4507
rect 13916 4489 13924 4499
rect 13869 4482 13924 4489
rect 13941 4482 13949 4499
rect 13869 4474 13949 4482
rect 14250 4483 14294 4491
rect 13869 4440 13884 4474
rect 14250 4466 14258 4483
rect 14275 4466 14294 4483
rect 14250 4458 14294 4466
rect 13905 4440 13920 4453
rect 14279 4440 14294 4458
rect 14315 4440 14330 4512
rect 14359 4440 14374 4564
rect 14403 4543 14418 4614
rect 14970 4597 14985 4614
rect 14960 4589 14993 4597
rect 14960 4572 14968 4589
rect 14985 4572 14993 4589
rect 14960 4564 14993 4572
rect 14395 4535 14428 4543
rect 14395 4518 14403 4535
rect 14420 4518 14428 4535
rect 14395 4510 14428 4518
rect 14861 4537 14894 4545
rect 14861 4520 14869 4537
rect 14886 4527 14894 4537
rect 14886 4520 14941 4527
rect 14861 4512 14941 4520
rect 14403 4440 14418 4510
rect 14494 4499 14527 4507
rect 14494 4489 14502 4499
rect 14447 4482 14502 4489
rect 14519 4482 14527 4499
rect 14447 4474 14527 4482
rect 14861 4483 14905 4491
rect 14447 4440 14462 4474
rect 14861 4466 14869 4483
rect 14886 4466 14905 4483
rect 14861 4458 14905 4466
rect 14483 4440 14498 4453
rect 14890 4440 14905 4458
rect 14926 4440 14941 4512
rect 14970 4440 14985 4564
rect 15014 4543 15029 4614
rect 15581 4597 15596 4614
rect 15571 4589 15604 4597
rect 15571 4572 15579 4589
rect 15596 4572 15604 4589
rect 15571 4564 15604 4572
rect 15006 4535 15039 4543
rect 15006 4518 15014 4535
rect 15031 4518 15039 4535
rect 15006 4510 15039 4518
rect 15472 4537 15505 4545
rect 15472 4520 15480 4537
rect 15497 4527 15505 4537
rect 15497 4520 15552 4527
rect 15472 4512 15552 4520
rect 15014 4440 15029 4510
rect 15105 4499 15138 4507
rect 15105 4489 15113 4499
rect 15058 4482 15113 4489
rect 15130 4482 15138 4499
rect 15058 4474 15138 4482
rect 15472 4483 15516 4491
rect 15058 4440 15073 4474
rect 15472 4466 15480 4483
rect 15497 4466 15516 4483
rect 15472 4458 15516 4466
rect 15094 4440 15109 4453
rect 15501 4440 15516 4458
rect 15537 4440 15552 4512
rect 15581 4440 15596 4564
rect 15625 4543 15640 4614
rect 15617 4535 15650 4543
rect 15617 4518 15625 4535
rect 15642 4518 15650 4535
rect 15617 4510 15650 4518
rect 15625 4440 15640 4510
rect 15716 4499 15749 4507
rect 15716 4489 15724 4499
rect 15669 4482 15724 4489
rect 15741 4482 15749 4499
rect 15669 4474 15749 4482
rect 15669 4440 15684 4474
rect 15705 4440 15720 4453
rect 12479 4306 12494 4340
rect 12515 4327 12530 4340
rect 12559 4327 12574 4340
rect 12603 4327 12618 4340
rect 12647 4327 12662 4340
rect 12683 4306 12698 4340
rect 12479 4291 12698 4306
rect 13090 4306 13105 4340
rect 13126 4327 13141 4340
rect 13170 4327 13185 4340
rect 13214 4327 13229 4340
rect 13258 4327 13273 4340
rect 13294 4306 13309 4340
rect 13090 4291 13309 4306
rect 13701 4306 13716 4340
rect 13737 4327 13752 4340
rect 13781 4327 13796 4340
rect 13825 4327 13840 4340
rect 13869 4327 13884 4340
rect 13905 4306 13920 4340
rect 13701 4291 13920 4306
rect 14279 4306 14294 4340
rect 14315 4327 14330 4340
rect 14359 4327 14374 4340
rect 14403 4327 14418 4340
rect 14447 4327 14462 4340
rect 14483 4306 14498 4340
rect 14279 4291 14498 4306
rect 14890 4306 14905 4340
rect 14926 4327 14941 4340
rect 14970 4327 14985 4340
rect 15014 4327 15029 4340
rect 15058 4327 15073 4340
rect 15094 4306 15109 4340
rect 14890 4291 15109 4306
rect 15501 4306 15516 4340
rect 15537 4327 15552 4340
rect 15581 4327 15596 4340
rect 15625 4327 15640 4340
rect 15669 4327 15684 4340
rect 15705 4306 15720 4340
rect 15501 4291 15720 4306
<< polycont >>
rect 13168 7802 13185 7819
rect 13069 7750 13086 7767
rect 13069 7696 13086 7713
rect 13779 7802 13796 7819
rect 13214 7748 13231 7765
rect 13680 7750 13697 7767
rect 13313 7712 13330 7729
rect 13680 7696 13697 7713
rect 14357 7802 14374 7819
rect 13825 7748 13842 7765
rect 14258 7750 14275 7767
rect 13924 7712 13941 7729
rect 14258 7696 14275 7713
rect 14968 7802 14985 7819
rect 14403 7748 14420 7765
rect 14869 7750 14886 7767
rect 14502 7712 14519 7729
rect 14869 7696 14886 7713
rect 15579 7802 15596 7819
rect 15014 7748 15031 7765
rect 15480 7750 15497 7767
rect 15113 7712 15130 7729
rect 15480 7696 15497 7713
rect 15625 7748 15642 7765
rect 15724 7712 15741 7729
rect 12557 7152 12574 7169
rect 12458 7100 12475 7117
rect 12458 7046 12475 7063
rect 13168 7152 13185 7169
rect 12603 7098 12620 7115
rect 13069 7100 13086 7117
rect 12702 7062 12719 7079
rect 13069 7046 13086 7063
rect 13779 7152 13796 7169
rect 13214 7098 13231 7115
rect 13680 7100 13697 7117
rect 13313 7062 13330 7079
rect 13680 7046 13697 7063
rect 14357 7152 14374 7169
rect 13825 7098 13842 7115
rect 14258 7100 14275 7117
rect 13924 7062 13941 7079
rect 14258 7046 14275 7063
rect 14968 7152 14985 7169
rect 14403 7098 14420 7115
rect 14869 7100 14886 7117
rect 14502 7062 14519 7079
rect 14869 7046 14886 7063
rect 15579 7152 15596 7169
rect 15014 7098 15031 7115
rect 15480 7100 15497 7117
rect 15113 7062 15130 7079
rect 15480 7046 15497 7063
rect 15625 7098 15642 7115
rect 15724 7062 15741 7079
rect 12557 6512 12574 6529
rect 12458 6460 12475 6477
rect 12458 6406 12475 6423
rect 13168 6512 13185 6529
rect 12603 6458 12620 6475
rect 13069 6460 13086 6477
rect 12702 6422 12719 6439
rect 13069 6406 13086 6423
rect 13779 6512 13796 6529
rect 13214 6458 13231 6475
rect 13680 6460 13697 6477
rect 13313 6422 13330 6439
rect 13680 6406 13697 6423
rect 14357 6512 14374 6529
rect 13825 6458 13842 6475
rect 14258 6460 14275 6477
rect 13924 6422 13941 6439
rect 14258 6406 14275 6423
rect 14968 6512 14985 6529
rect 14403 6458 14420 6475
rect 14869 6460 14886 6477
rect 14502 6422 14519 6439
rect 14869 6406 14886 6423
rect 15579 6512 15596 6529
rect 15014 6458 15031 6475
rect 15480 6460 15497 6477
rect 15113 6422 15130 6439
rect 15480 6406 15497 6423
rect 15625 6458 15642 6475
rect 15724 6422 15741 6439
rect 12557 5862 12574 5879
rect 12458 5810 12475 5827
rect 12458 5756 12475 5773
rect 13168 5862 13185 5879
rect 12603 5808 12620 5825
rect 13069 5810 13086 5827
rect 12702 5772 12719 5789
rect 13069 5756 13086 5773
rect 13779 5862 13796 5879
rect 13214 5808 13231 5825
rect 13680 5810 13697 5827
rect 13313 5772 13330 5789
rect 13680 5756 13697 5773
rect 14357 5862 14374 5879
rect 13825 5808 13842 5825
rect 14258 5810 14275 5827
rect 13924 5772 13941 5789
rect 14258 5756 14275 5773
rect 14968 5862 14985 5879
rect 14403 5808 14420 5825
rect 14869 5810 14886 5827
rect 14502 5772 14519 5789
rect 14869 5756 14886 5773
rect 15579 5862 15596 5879
rect 15014 5808 15031 5825
rect 15480 5810 15497 5827
rect 15113 5772 15130 5789
rect 15480 5756 15497 5773
rect 15625 5808 15642 5825
rect 15724 5772 15741 5789
rect 12557 5212 12574 5229
rect 12458 5160 12475 5177
rect 12458 5106 12475 5123
rect 13168 5212 13185 5229
rect 12603 5158 12620 5175
rect 13069 5160 13086 5177
rect 12702 5122 12719 5139
rect 13069 5106 13086 5123
rect 13779 5212 13796 5229
rect 13214 5158 13231 5175
rect 13680 5160 13697 5177
rect 13313 5122 13330 5139
rect 13680 5106 13697 5123
rect 14357 5212 14374 5229
rect 13825 5158 13842 5175
rect 14258 5160 14275 5177
rect 13924 5122 13941 5139
rect 14258 5106 14275 5123
rect 14968 5212 14985 5229
rect 14403 5158 14420 5175
rect 14869 5160 14886 5177
rect 14502 5122 14519 5139
rect 14869 5106 14886 5123
rect 15579 5212 15596 5229
rect 15014 5158 15031 5175
rect 15480 5160 15497 5177
rect 15113 5122 15130 5139
rect 15480 5106 15497 5123
rect 15625 5158 15642 5175
rect 15724 5122 15741 5139
rect 12557 4572 12574 4589
rect 12458 4520 12475 4537
rect 12458 4466 12475 4483
rect 13168 4572 13185 4589
rect 12603 4518 12620 4535
rect 13069 4520 13086 4537
rect 12702 4482 12719 4499
rect 13069 4466 13086 4483
rect 13779 4572 13796 4589
rect 13214 4518 13231 4535
rect 13680 4520 13697 4537
rect 13313 4482 13330 4499
rect 13680 4466 13697 4483
rect 14357 4572 14374 4589
rect 13825 4518 13842 4535
rect 14258 4520 14275 4537
rect 13924 4482 13941 4499
rect 14258 4466 14275 4483
rect 14968 4572 14985 4589
rect 14403 4518 14420 4535
rect 14869 4520 14886 4537
rect 14502 4482 14519 4499
rect 14869 4466 14886 4483
rect 15579 4572 15596 4589
rect 15014 4518 15031 4535
rect 15480 4520 15497 4537
rect 15113 4482 15130 4499
rect 15480 4466 15497 4483
rect 15625 4518 15642 4535
rect 15724 4482 15741 4499
<< locali >>
rect 13186 8062 13190 8081
rect 13209 8062 13213 8081
rect 13111 8039 13169 8047
rect 13111 8022 13147 8039
rect 13164 8022 13169 8039
rect 13111 8005 13169 8022
rect 13111 7988 13147 8005
rect 13164 7988 13169 8005
rect 13111 7971 13169 7988
rect 13111 7954 13147 7971
rect 13164 7954 13169 7971
rect 13111 7937 13169 7954
rect 13111 7920 13147 7937
rect 13164 7920 13169 7937
rect 13111 7903 13169 7920
rect 13111 7886 13147 7903
rect 13164 7886 13169 7903
rect 13111 7869 13169 7886
rect 13111 7852 13147 7869
rect 13164 7852 13169 7869
rect 13111 7844 13169 7852
rect 13186 8039 13213 8062
rect 13797 8062 13801 8081
rect 13820 8062 13824 8081
rect 13186 8022 13191 8039
rect 13208 8022 13213 8039
rect 13186 8005 13213 8022
rect 13186 7988 13191 8005
rect 13208 7988 13213 8005
rect 13186 7971 13213 7988
rect 13186 7954 13191 7971
rect 13208 7954 13213 7971
rect 13186 7937 13213 7954
rect 13186 7920 13191 7937
rect 13208 7920 13213 7937
rect 13186 7903 13213 7920
rect 13186 7886 13191 7903
rect 13208 7886 13213 7903
rect 13186 7869 13213 7886
rect 13186 7852 13191 7869
rect 13208 7852 13213 7869
rect 13186 7844 13213 7852
rect 13230 8039 13288 8047
rect 13230 8022 13235 8039
rect 13252 8022 13288 8039
rect 13230 8005 13288 8022
rect 13230 7988 13235 8005
rect 13252 7988 13288 8005
rect 13230 7971 13288 7988
rect 13230 7954 13235 7971
rect 13252 7954 13288 7971
rect 13230 7937 13288 7954
rect 13230 7920 13235 7937
rect 13252 7920 13288 7937
rect 13230 7903 13288 7920
rect 13230 7886 13235 7903
rect 13252 7886 13288 7903
rect 13230 7869 13288 7886
rect 13230 7852 13235 7869
rect 13252 7852 13288 7869
rect 13230 7844 13288 7852
rect 13061 7767 13094 7775
rect 13061 7750 13069 7767
rect 13086 7750 13094 7767
rect 13061 7742 13094 7750
rect 13111 7757 13138 7844
rect 13160 7819 13193 7827
rect 13160 7802 13168 7819
rect 13185 7811 13193 7819
rect 13261 7811 13288 7844
rect 13185 7802 13288 7811
rect 13160 7794 13288 7802
rect 13206 7765 13239 7773
rect 13206 7757 13214 7765
rect 13111 7748 13214 7757
rect 13231 7748 13239 7765
rect 13111 7740 13239 7748
rect 13061 7713 13094 7721
rect 13061 7696 13069 7713
rect 13086 7696 13094 7713
rect 13061 7688 13094 7696
rect 13111 7671 13138 7740
rect 13261 7671 13288 7794
rect 13722 8039 13780 8047
rect 13722 8022 13758 8039
rect 13775 8022 13780 8039
rect 13722 8005 13780 8022
rect 13722 7988 13758 8005
rect 13775 7988 13780 8005
rect 13722 7971 13780 7988
rect 13722 7954 13758 7971
rect 13775 7954 13780 7971
rect 13722 7937 13780 7954
rect 13722 7920 13758 7937
rect 13775 7920 13780 7937
rect 13722 7903 13780 7920
rect 13722 7886 13758 7903
rect 13775 7886 13780 7903
rect 13722 7869 13780 7886
rect 13722 7852 13758 7869
rect 13775 7852 13780 7869
rect 13722 7844 13780 7852
rect 13797 8039 13824 8062
rect 14375 8062 14379 8081
rect 14398 8062 14402 8081
rect 13797 8022 13802 8039
rect 13819 8022 13824 8039
rect 13797 8005 13824 8022
rect 13797 7988 13802 8005
rect 13819 7988 13824 8005
rect 13797 7971 13824 7988
rect 13797 7954 13802 7971
rect 13819 7954 13824 7971
rect 13797 7937 13824 7954
rect 13797 7920 13802 7937
rect 13819 7920 13824 7937
rect 13797 7903 13824 7920
rect 13797 7886 13802 7903
rect 13819 7886 13824 7903
rect 13797 7869 13824 7886
rect 13797 7852 13802 7869
rect 13819 7852 13824 7869
rect 13797 7844 13824 7852
rect 13841 8039 13899 8047
rect 13841 8022 13846 8039
rect 13863 8022 13899 8039
rect 13841 8005 13899 8022
rect 13841 7988 13846 8005
rect 13863 7988 13899 8005
rect 13841 7971 13899 7988
rect 13841 7954 13846 7971
rect 13863 7954 13899 7971
rect 13841 7937 13899 7954
rect 13841 7920 13846 7937
rect 13863 7920 13899 7937
rect 13841 7903 13899 7920
rect 13841 7886 13846 7903
rect 13863 7886 13899 7903
rect 13841 7869 13899 7886
rect 13841 7852 13846 7869
rect 13863 7852 13899 7869
rect 13841 7844 13899 7852
rect 13672 7767 13705 7775
rect 13672 7750 13680 7767
rect 13697 7750 13705 7767
rect 13672 7742 13705 7750
rect 13722 7757 13749 7844
rect 13771 7819 13804 7827
rect 13771 7802 13779 7819
rect 13796 7811 13804 7819
rect 13872 7811 13899 7844
rect 13796 7802 13899 7811
rect 13771 7794 13899 7802
rect 13817 7765 13850 7773
rect 13817 7757 13825 7765
rect 13722 7748 13825 7757
rect 13842 7748 13850 7765
rect 13722 7740 13850 7748
rect 13305 7729 13338 7737
rect 13305 7712 13313 7729
rect 13330 7712 13338 7729
rect 13305 7704 13338 7712
rect 13672 7713 13705 7721
rect 13672 7696 13680 7713
rect 13697 7696 13705 7713
rect 13672 7688 13705 7696
rect 13722 7671 13749 7740
rect 13872 7671 13899 7794
rect 14300 8039 14358 8047
rect 14300 8022 14336 8039
rect 14353 8022 14358 8039
rect 14300 8005 14358 8022
rect 14300 7988 14336 8005
rect 14353 7988 14358 8005
rect 14300 7971 14358 7988
rect 14300 7954 14336 7971
rect 14353 7954 14358 7971
rect 14300 7937 14358 7954
rect 14300 7920 14336 7937
rect 14353 7920 14358 7937
rect 14300 7903 14358 7920
rect 14300 7886 14336 7903
rect 14353 7886 14358 7903
rect 14300 7869 14358 7886
rect 14300 7852 14336 7869
rect 14353 7852 14358 7869
rect 14300 7844 14358 7852
rect 14375 8039 14402 8062
rect 14986 8062 14990 8081
rect 15009 8062 15013 8081
rect 14375 8022 14380 8039
rect 14397 8022 14402 8039
rect 14375 8005 14402 8022
rect 14375 7988 14380 8005
rect 14397 7988 14402 8005
rect 14375 7971 14402 7988
rect 14375 7954 14380 7971
rect 14397 7954 14402 7971
rect 14375 7937 14402 7954
rect 14375 7920 14380 7937
rect 14397 7920 14402 7937
rect 14375 7903 14402 7920
rect 14375 7886 14380 7903
rect 14397 7886 14402 7903
rect 14375 7869 14402 7886
rect 14375 7852 14380 7869
rect 14397 7852 14402 7869
rect 14375 7844 14402 7852
rect 14419 8039 14477 8047
rect 14419 8022 14424 8039
rect 14441 8022 14477 8039
rect 14419 8005 14477 8022
rect 14419 7988 14424 8005
rect 14441 7988 14477 8005
rect 14419 7971 14477 7988
rect 14419 7954 14424 7971
rect 14441 7954 14477 7971
rect 14419 7937 14477 7954
rect 14419 7920 14424 7937
rect 14441 7920 14477 7937
rect 14419 7903 14477 7920
rect 14419 7886 14424 7903
rect 14441 7886 14477 7903
rect 14419 7869 14477 7886
rect 14419 7852 14424 7869
rect 14441 7852 14477 7869
rect 14419 7844 14477 7852
rect 14250 7767 14283 7775
rect 14250 7750 14258 7767
rect 14275 7750 14283 7767
rect 14250 7742 14283 7750
rect 14300 7757 14327 7844
rect 14349 7819 14382 7827
rect 14349 7802 14357 7819
rect 14374 7811 14382 7819
rect 14450 7811 14477 7844
rect 14374 7802 14477 7811
rect 14349 7794 14477 7802
rect 14395 7765 14428 7773
rect 14395 7757 14403 7765
rect 14300 7748 14403 7757
rect 14420 7748 14428 7765
rect 14300 7740 14428 7748
rect 13916 7729 13949 7737
rect 13916 7712 13924 7729
rect 13941 7712 13949 7729
rect 13916 7704 13949 7712
rect 14250 7713 14283 7721
rect 14250 7696 14258 7713
rect 14275 7696 14283 7713
rect 14250 7688 14283 7696
rect 14300 7671 14327 7740
rect 14450 7671 14477 7794
rect 14911 8039 14969 8047
rect 14911 8022 14947 8039
rect 14964 8022 14969 8039
rect 14911 8005 14969 8022
rect 14911 7988 14947 8005
rect 14964 7988 14969 8005
rect 14911 7971 14969 7988
rect 14911 7954 14947 7971
rect 14964 7954 14969 7971
rect 14911 7937 14969 7954
rect 14911 7920 14947 7937
rect 14964 7920 14969 7937
rect 14911 7903 14969 7920
rect 14911 7886 14947 7903
rect 14964 7886 14969 7903
rect 14911 7869 14969 7886
rect 14911 7852 14947 7869
rect 14964 7852 14969 7869
rect 14911 7844 14969 7852
rect 14986 8039 15013 8062
rect 15597 8062 15601 8081
rect 15620 8062 15624 8081
rect 14986 8022 14991 8039
rect 15008 8022 15013 8039
rect 14986 8005 15013 8022
rect 14986 7988 14991 8005
rect 15008 7988 15013 8005
rect 14986 7971 15013 7988
rect 14986 7954 14991 7971
rect 15008 7954 15013 7971
rect 14986 7937 15013 7954
rect 14986 7920 14991 7937
rect 15008 7920 15013 7937
rect 14986 7903 15013 7920
rect 14986 7886 14991 7903
rect 15008 7886 15013 7903
rect 14986 7869 15013 7886
rect 14986 7852 14991 7869
rect 15008 7852 15013 7869
rect 14986 7844 15013 7852
rect 15030 8039 15088 8047
rect 15030 8022 15035 8039
rect 15052 8022 15088 8039
rect 15030 8005 15088 8022
rect 15030 7988 15035 8005
rect 15052 7988 15088 8005
rect 15030 7971 15088 7988
rect 15030 7954 15035 7971
rect 15052 7954 15088 7971
rect 15030 7937 15088 7954
rect 15030 7920 15035 7937
rect 15052 7920 15088 7937
rect 15030 7903 15088 7920
rect 15030 7886 15035 7903
rect 15052 7886 15088 7903
rect 15030 7869 15088 7886
rect 15030 7852 15035 7869
rect 15052 7852 15088 7869
rect 15030 7844 15088 7852
rect 14861 7767 14894 7775
rect 14861 7750 14869 7767
rect 14886 7750 14894 7767
rect 14861 7742 14894 7750
rect 14911 7757 14938 7844
rect 14960 7819 14993 7827
rect 14960 7802 14968 7819
rect 14985 7811 14993 7819
rect 15061 7811 15088 7844
rect 14985 7802 15088 7811
rect 14960 7794 15088 7802
rect 15006 7765 15039 7773
rect 15006 7757 15014 7765
rect 14911 7748 15014 7757
rect 15031 7748 15039 7765
rect 14911 7740 15039 7748
rect 14494 7729 14527 7737
rect 14494 7712 14502 7729
rect 14519 7712 14527 7729
rect 14494 7704 14527 7712
rect 14861 7713 14894 7721
rect 14861 7696 14869 7713
rect 14886 7696 14894 7713
rect 14861 7688 14894 7696
rect 14911 7671 14938 7740
rect 15061 7671 15088 7794
rect 15522 8039 15580 8047
rect 15522 8022 15558 8039
rect 15575 8022 15580 8039
rect 15522 8005 15580 8022
rect 15522 7988 15558 8005
rect 15575 7988 15580 8005
rect 15522 7971 15580 7988
rect 15522 7954 15558 7971
rect 15575 7954 15580 7971
rect 15522 7937 15580 7954
rect 15522 7920 15558 7937
rect 15575 7920 15580 7937
rect 15522 7903 15580 7920
rect 15522 7886 15558 7903
rect 15575 7886 15580 7903
rect 15522 7869 15580 7886
rect 15522 7852 15558 7869
rect 15575 7852 15580 7869
rect 15522 7844 15580 7852
rect 15597 8039 15624 8062
rect 15597 8022 15602 8039
rect 15619 8022 15624 8039
rect 15597 8005 15624 8022
rect 15597 7988 15602 8005
rect 15619 7988 15624 8005
rect 15597 7971 15624 7988
rect 15597 7954 15602 7971
rect 15619 7954 15624 7971
rect 15597 7937 15624 7954
rect 15597 7920 15602 7937
rect 15619 7920 15624 7937
rect 15597 7903 15624 7920
rect 15597 7886 15602 7903
rect 15619 7886 15624 7903
rect 15597 7869 15624 7886
rect 15597 7852 15602 7869
rect 15619 7852 15624 7869
rect 15597 7844 15624 7852
rect 15641 8039 15699 8047
rect 15641 8022 15646 8039
rect 15663 8022 15699 8039
rect 15641 8005 15699 8022
rect 15641 7988 15646 8005
rect 15663 7988 15699 8005
rect 15641 7971 15699 7988
rect 15641 7954 15646 7971
rect 15663 7954 15699 7971
rect 15641 7937 15699 7954
rect 15641 7920 15646 7937
rect 15663 7920 15699 7937
rect 15641 7903 15699 7920
rect 15641 7886 15646 7903
rect 15663 7886 15699 7903
rect 15641 7869 15699 7886
rect 15641 7852 15646 7869
rect 15663 7852 15699 7869
rect 15641 7844 15699 7852
rect 15472 7767 15505 7775
rect 15472 7750 15480 7767
rect 15497 7750 15505 7767
rect 15472 7742 15505 7750
rect 15522 7757 15549 7844
rect 15571 7819 15604 7827
rect 15571 7802 15579 7819
rect 15596 7811 15604 7819
rect 15672 7811 15699 7844
rect 15596 7802 15699 7811
rect 15571 7794 15699 7802
rect 15617 7765 15650 7773
rect 15617 7757 15625 7765
rect 15522 7748 15625 7757
rect 15642 7748 15650 7765
rect 15522 7740 15650 7748
rect 15105 7729 15138 7737
rect 15105 7712 15113 7729
rect 15130 7712 15138 7729
rect 15105 7704 15138 7712
rect 15472 7713 15505 7721
rect 15472 7696 15480 7713
rect 15497 7696 15505 7713
rect 15472 7688 15505 7696
rect 15522 7671 15549 7740
rect 15672 7671 15699 7794
rect 15716 7729 15749 7737
rect 15716 7712 15724 7729
rect 15741 7712 15749 7729
rect 15716 7704 15749 7712
rect 13062 7663 13089 7671
rect 13062 7646 13067 7663
rect 13084 7646 13089 7663
rect 13062 7629 13089 7646
rect 13062 7612 13067 7629
rect 13084 7612 13089 7629
rect 13062 7595 13089 7612
rect 13062 7578 13067 7595
rect 13084 7578 13089 7595
rect 13062 7570 13089 7578
rect 13111 7663 13169 7671
rect 13111 7646 13147 7663
rect 13164 7646 13169 7663
rect 13111 7629 13169 7646
rect 13111 7612 13147 7629
rect 13164 7612 13169 7629
rect 13111 7595 13169 7612
rect 13111 7578 13147 7595
rect 13164 7578 13169 7595
rect 13111 7570 13169 7578
rect 13186 7663 13213 7671
rect 13186 7646 13191 7663
rect 13208 7646 13213 7663
rect 13186 7629 13213 7646
rect 13186 7612 13191 7629
rect 13208 7612 13213 7629
rect 13186 7595 13213 7612
rect 13186 7578 13191 7595
rect 13208 7578 13213 7595
rect 13186 7555 13213 7578
rect 13230 7663 13288 7671
rect 13230 7646 13235 7663
rect 13252 7646 13288 7663
rect 13230 7629 13288 7646
rect 13230 7612 13235 7629
rect 13252 7612 13288 7629
rect 13230 7595 13288 7612
rect 13230 7578 13235 7595
rect 13252 7578 13288 7595
rect 13230 7570 13288 7578
rect 13310 7663 13337 7671
rect 13310 7646 13315 7663
rect 13332 7646 13337 7663
rect 13310 7629 13337 7646
rect 13310 7612 13315 7629
rect 13332 7612 13337 7629
rect 13310 7595 13337 7612
rect 13310 7578 13315 7595
rect 13332 7578 13337 7595
rect 13310 7570 13337 7578
rect 13673 7663 13700 7671
rect 13673 7646 13678 7663
rect 13695 7646 13700 7663
rect 13673 7629 13700 7646
rect 13673 7612 13678 7629
rect 13695 7612 13700 7629
rect 13673 7595 13700 7612
rect 13673 7578 13678 7595
rect 13695 7578 13700 7595
rect 13673 7570 13700 7578
rect 13722 7663 13780 7671
rect 13722 7646 13758 7663
rect 13775 7646 13780 7663
rect 13722 7629 13780 7646
rect 13722 7612 13758 7629
rect 13775 7612 13780 7629
rect 13722 7595 13780 7612
rect 13722 7578 13758 7595
rect 13775 7578 13780 7595
rect 13722 7570 13780 7578
rect 13797 7663 13824 7671
rect 13797 7646 13802 7663
rect 13819 7646 13824 7663
rect 13797 7629 13824 7646
rect 13797 7612 13802 7629
rect 13819 7612 13824 7629
rect 13797 7595 13824 7612
rect 13797 7578 13802 7595
rect 13819 7578 13824 7595
rect 13186 7536 13190 7555
rect 13209 7536 13213 7555
rect 13797 7555 13824 7578
rect 13841 7663 13899 7671
rect 13841 7646 13846 7663
rect 13863 7646 13899 7663
rect 13841 7629 13899 7646
rect 13841 7612 13846 7629
rect 13863 7612 13899 7629
rect 13841 7595 13899 7612
rect 13841 7578 13846 7595
rect 13863 7578 13899 7595
rect 13841 7570 13899 7578
rect 13921 7663 13948 7671
rect 13921 7646 13926 7663
rect 13943 7646 13948 7663
rect 13921 7629 13948 7646
rect 13921 7612 13926 7629
rect 13943 7612 13948 7629
rect 13921 7595 13948 7612
rect 13921 7578 13926 7595
rect 13943 7578 13948 7595
rect 13921 7570 13948 7578
rect 14251 7663 14278 7671
rect 14251 7646 14256 7663
rect 14273 7646 14278 7663
rect 14251 7629 14278 7646
rect 14251 7612 14256 7629
rect 14273 7612 14278 7629
rect 14251 7595 14278 7612
rect 14251 7578 14256 7595
rect 14273 7578 14278 7595
rect 14251 7570 14278 7578
rect 14300 7663 14358 7671
rect 14300 7646 14336 7663
rect 14353 7646 14358 7663
rect 14300 7629 14358 7646
rect 14300 7612 14336 7629
rect 14353 7612 14358 7629
rect 14300 7595 14358 7612
rect 14300 7578 14336 7595
rect 14353 7578 14358 7595
rect 14300 7570 14358 7578
rect 14375 7663 14402 7671
rect 14375 7646 14380 7663
rect 14397 7646 14402 7663
rect 14375 7629 14402 7646
rect 14375 7612 14380 7629
rect 14397 7612 14402 7629
rect 14375 7595 14402 7612
rect 14375 7578 14380 7595
rect 14397 7578 14402 7595
rect 13797 7536 13801 7555
rect 13820 7536 13824 7555
rect 14375 7555 14402 7578
rect 14419 7663 14477 7671
rect 14419 7646 14424 7663
rect 14441 7646 14477 7663
rect 14419 7629 14477 7646
rect 14419 7612 14424 7629
rect 14441 7612 14477 7629
rect 14419 7595 14477 7612
rect 14419 7578 14424 7595
rect 14441 7578 14477 7595
rect 14419 7570 14477 7578
rect 14499 7663 14526 7671
rect 14499 7646 14504 7663
rect 14521 7646 14526 7663
rect 14499 7629 14526 7646
rect 14499 7612 14504 7629
rect 14521 7612 14526 7629
rect 14499 7595 14526 7612
rect 14499 7578 14504 7595
rect 14521 7578 14526 7595
rect 14499 7570 14526 7578
rect 14862 7663 14889 7671
rect 14862 7646 14867 7663
rect 14884 7646 14889 7663
rect 14862 7629 14889 7646
rect 14862 7612 14867 7629
rect 14884 7612 14889 7629
rect 14862 7595 14889 7612
rect 14862 7578 14867 7595
rect 14884 7578 14889 7595
rect 14862 7570 14889 7578
rect 14911 7663 14969 7671
rect 14911 7646 14947 7663
rect 14964 7646 14969 7663
rect 14911 7629 14969 7646
rect 14911 7612 14947 7629
rect 14964 7612 14969 7629
rect 14911 7595 14969 7612
rect 14911 7578 14947 7595
rect 14964 7578 14969 7595
rect 14911 7570 14969 7578
rect 14986 7663 15013 7671
rect 14986 7646 14991 7663
rect 15008 7646 15013 7663
rect 14986 7629 15013 7646
rect 14986 7612 14991 7629
rect 15008 7612 15013 7629
rect 14986 7595 15013 7612
rect 14986 7578 14991 7595
rect 15008 7578 15013 7595
rect 14375 7536 14379 7555
rect 14398 7536 14402 7555
rect 14986 7555 15013 7578
rect 15030 7663 15088 7671
rect 15030 7646 15035 7663
rect 15052 7646 15088 7663
rect 15030 7629 15088 7646
rect 15030 7612 15035 7629
rect 15052 7612 15088 7629
rect 15030 7595 15088 7612
rect 15030 7578 15035 7595
rect 15052 7578 15088 7595
rect 15030 7570 15088 7578
rect 15110 7663 15137 7671
rect 15110 7646 15115 7663
rect 15132 7646 15137 7663
rect 15110 7629 15137 7646
rect 15110 7612 15115 7629
rect 15132 7612 15137 7629
rect 15110 7595 15137 7612
rect 15110 7578 15115 7595
rect 15132 7578 15137 7595
rect 15110 7570 15137 7578
rect 15473 7663 15500 7671
rect 15473 7646 15478 7663
rect 15495 7646 15500 7663
rect 15473 7629 15500 7646
rect 15473 7612 15478 7629
rect 15495 7612 15500 7629
rect 15473 7595 15500 7612
rect 15473 7578 15478 7595
rect 15495 7578 15500 7595
rect 15473 7570 15500 7578
rect 15522 7663 15580 7671
rect 15522 7646 15558 7663
rect 15575 7646 15580 7663
rect 15522 7629 15580 7646
rect 15522 7612 15558 7629
rect 15575 7612 15580 7629
rect 15522 7595 15580 7612
rect 15522 7578 15558 7595
rect 15575 7578 15580 7595
rect 15522 7570 15580 7578
rect 15597 7663 15624 7671
rect 15597 7646 15602 7663
rect 15619 7646 15624 7663
rect 15597 7629 15624 7646
rect 15597 7612 15602 7629
rect 15619 7612 15624 7629
rect 15597 7595 15624 7612
rect 15597 7578 15602 7595
rect 15619 7578 15624 7595
rect 14986 7536 14990 7555
rect 15009 7536 15013 7555
rect 15597 7555 15624 7578
rect 15641 7663 15699 7671
rect 15641 7646 15646 7663
rect 15663 7646 15699 7663
rect 15641 7629 15699 7646
rect 15641 7612 15646 7629
rect 15663 7612 15699 7629
rect 15641 7595 15699 7612
rect 15641 7578 15646 7595
rect 15663 7578 15699 7595
rect 15641 7570 15699 7578
rect 15721 7663 15748 7671
rect 15721 7646 15726 7663
rect 15743 7646 15748 7663
rect 15721 7629 15748 7646
rect 15721 7612 15726 7629
rect 15743 7612 15748 7629
rect 15721 7595 15748 7612
rect 15721 7578 15726 7595
rect 15743 7578 15748 7595
rect 15721 7570 15748 7578
rect 15597 7536 15601 7555
rect 15620 7536 15624 7555
rect 12575 7412 12579 7431
rect 12598 7412 12602 7431
rect 12500 7389 12558 7397
rect 12500 7372 12536 7389
rect 12553 7372 12558 7389
rect 12500 7355 12558 7372
rect 12500 7338 12536 7355
rect 12553 7338 12558 7355
rect 12500 7321 12558 7338
rect 12500 7304 12536 7321
rect 12553 7304 12558 7321
rect 12500 7287 12558 7304
rect 12500 7270 12536 7287
rect 12553 7270 12558 7287
rect 12500 7253 12558 7270
rect 12500 7236 12536 7253
rect 12553 7236 12558 7253
rect 12500 7219 12558 7236
rect 12500 7202 12536 7219
rect 12553 7202 12558 7219
rect 12500 7194 12558 7202
rect 12575 7389 12602 7412
rect 13186 7412 13190 7431
rect 13209 7412 13213 7431
rect 12575 7372 12580 7389
rect 12597 7372 12602 7389
rect 12575 7355 12602 7372
rect 12575 7338 12580 7355
rect 12597 7338 12602 7355
rect 12575 7321 12602 7338
rect 12575 7304 12580 7321
rect 12597 7304 12602 7321
rect 12575 7287 12602 7304
rect 12575 7270 12580 7287
rect 12597 7270 12602 7287
rect 12575 7253 12602 7270
rect 12575 7236 12580 7253
rect 12597 7236 12602 7253
rect 12575 7219 12602 7236
rect 12575 7202 12580 7219
rect 12597 7202 12602 7219
rect 12575 7194 12602 7202
rect 12619 7389 12677 7397
rect 12619 7372 12624 7389
rect 12641 7372 12677 7389
rect 12619 7355 12677 7372
rect 12619 7338 12624 7355
rect 12641 7338 12677 7355
rect 12619 7321 12677 7338
rect 12619 7304 12624 7321
rect 12641 7304 12677 7321
rect 12619 7287 12677 7304
rect 12619 7270 12624 7287
rect 12641 7270 12677 7287
rect 12619 7253 12677 7270
rect 12619 7236 12624 7253
rect 12641 7236 12677 7253
rect 12619 7219 12677 7236
rect 12619 7202 12624 7219
rect 12641 7202 12677 7219
rect 12619 7194 12677 7202
rect 12450 7117 12483 7125
rect 12450 7100 12458 7117
rect 12475 7100 12483 7117
rect 12450 7092 12483 7100
rect 12500 7107 12527 7194
rect 12549 7169 12582 7177
rect 12549 7152 12557 7169
rect 12574 7161 12582 7169
rect 12650 7161 12677 7194
rect 12574 7152 12677 7161
rect 12549 7144 12677 7152
rect 12595 7115 12628 7123
rect 12595 7107 12603 7115
rect 12500 7098 12603 7107
rect 12620 7098 12628 7115
rect 12500 7090 12628 7098
rect 12450 7063 12483 7071
rect 12450 7046 12458 7063
rect 12475 7046 12483 7063
rect 12450 7038 12483 7046
rect 12500 7021 12527 7090
rect 12650 7021 12677 7144
rect 13111 7389 13169 7397
rect 13111 7372 13147 7389
rect 13164 7372 13169 7389
rect 13111 7355 13169 7372
rect 13111 7338 13147 7355
rect 13164 7338 13169 7355
rect 13111 7321 13169 7338
rect 13111 7304 13147 7321
rect 13164 7304 13169 7321
rect 13111 7287 13169 7304
rect 13111 7270 13147 7287
rect 13164 7270 13169 7287
rect 13111 7253 13169 7270
rect 13111 7236 13147 7253
rect 13164 7236 13169 7253
rect 13111 7219 13169 7236
rect 13111 7202 13147 7219
rect 13164 7202 13169 7219
rect 13111 7194 13169 7202
rect 13186 7389 13213 7412
rect 13797 7412 13801 7431
rect 13820 7412 13824 7431
rect 13186 7372 13191 7389
rect 13208 7372 13213 7389
rect 13186 7355 13213 7372
rect 13186 7338 13191 7355
rect 13208 7338 13213 7355
rect 13186 7321 13213 7338
rect 13186 7304 13191 7321
rect 13208 7304 13213 7321
rect 13186 7287 13213 7304
rect 13186 7270 13191 7287
rect 13208 7270 13213 7287
rect 13186 7253 13213 7270
rect 13186 7236 13191 7253
rect 13208 7236 13213 7253
rect 13186 7219 13213 7236
rect 13186 7202 13191 7219
rect 13208 7202 13213 7219
rect 13186 7194 13213 7202
rect 13230 7389 13288 7397
rect 13230 7372 13235 7389
rect 13252 7372 13288 7389
rect 13230 7355 13288 7372
rect 13230 7338 13235 7355
rect 13252 7338 13288 7355
rect 13230 7321 13288 7338
rect 13230 7304 13235 7321
rect 13252 7304 13288 7321
rect 13230 7287 13288 7304
rect 13230 7270 13235 7287
rect 13252 7270 13288 7287
rect 13230 7253 13288 7270
rect 13230 7236 13235 7253
rect 13252 7236 13288 7253
rect 13230 7219 13288 7236
rect 13230 7202 13235 7219
rect 13252 7202 13288 7219
rect 13230 7194 13288 7202
rect 13061 7117 13094 7125
rect 13061 7100 13069 7117
rect 13086 7100 13094 7117
rect 13061 7092 13094 7100
rect 13111 7107 13138 7194
rect 13160 7169 13193 7177
rect 13160 7152 13168 7169
rect 13185 7161 13193 7169
rect 13261 7161 13288 7194
rect 13185 7152 13288 7161
rect 13160 7144 13288 7152
rect 13206 7115 13239 7123
rect 13206 7107 13214 7115
rect 13111 7098 13214 7107
rect 13231 7098 13239 7115
rect 13111 7090 13239 7098
rect 12694 7079 12727 7087
rect 12694 7062 12702 7079
rect 12719 7062 12727 7079
rect 12694 7054 12727 7062
rect 13061 7063 13094 7071
rect 13061 7046 13069 7063
rect 13086 7046 13094 7063
rect 13061 7038 13094 7046
rect 13111 7021 13138 7090
rect 13261 7021 13288 7144
rect 13722 7389 13780 7397
rect 13722 7372 13758 7389
rect 13775 7372 13780 7389
rect 13722 7355 13780 7372
rect 13722 7338 13758 7355
rect 13775 7338 13780 7355
rect 13722 7321 13780 7338
rect 13722 7304 13758 7321
rect 13775 7304 13780 7321
rect 13722 7287 13780 7304
rect 13722 7270 13758 7287
rect 13775 7270 13780 7287
rect 13722 7253 13780 7270
rect 13722 7236 13758 7253
rect 13775 7236 13780 7253
rect 13722 7219 13780 7236
rect 13722 7202 13758 7219
rect 13775 7202 13780 7219
rect 13722 7194 13780 7202
rect 13797 7389 13824 7412
rect 14375 7412 14379 7431
rect 14398 7412 14402 7431
rect 13797 7372 13802 7389
rect 13819 7372 13824 7389
rect 13797 7355 13824 7372
rect 13797 7338 13802 7355
rect 13819 7338 13824 7355
rect 13797 7321 13824 7338
rect 13797 7304 13802 7321
rect 13819 7304 13824 7321
rect 13797 7287 13824 7304
rect 13797 7270 13802 7287
rect 13819 7270 13824 7287
rect 13797 7253 13824 7270
rect 13797 7236 13802 7253
rect 13819 7236 13824 7253
rect 13797 7219 13824 7236
rect 13797 7202 13802 7219
rect 13819 7202 13824 7219
rect 13797 7194 13824 7202
rect 13841 7389 13899 7397
rect 13841 7372 13846 7389
rect 13863 7372 13899 7389
rect 13841 7355 13899 7372
rect 13841 7338 13846 7355
rect 13863 7338 13899 7355
rect 13841 7321 13899 7338
rect 13841 7304 13846 7321
rect 13863 7304 13899 7321
rect 13841 7287 13899 7304
rect 13841 7270 13846 7287
rect 13863 7270 13899 7287
rect 13841 7253 13899 7270
rect 13841 7236 13846 7253
rect 13863 7236 13899 7253
rect 13841 7219 13899 7236
rect 13841 7202 13846 7219
rect 13863 7202 13899 7219
rect 13841 7194 13899 7202
rect 13672 7117 13705 7125
rect 13672 7100 13680 7117
rect 13697 7100 13705 7117
rect 13672 7092 13705 7100
rect 13722 7107 13749 7194
rect 13771 7169 13804 7177
rect 13771 7152 13779 7169
rect 13796 7161 13804 7169
rect 13872 7161 13899 7194
rect 13796 7152 13899 7161
rect 13771 7144 13899 7152
rect 13817 7115 13850 7123
rect 13817 7107 13825 7115
rect 13722 7098 13825 7107
rect 13842 7098 13850 7115
rect 13722 7090 13850 7098
rect 13305 7079 13338 7087
rect 13305 7062 13313 7079
rect 13330 7062 13338 7079
rect 13305 7054 13338 7062
rect 13672 7063 13705 7071
rect 13672 7046 13680 7063
rect 13697 7046 13705 7063
rect 13672 7038 13705 7046
rect 13722 7021 13749 7090
rect 13872 7021 13899 7144
rect 14300 7389 14358 7397
rect 14300 7372 14336 7389
rect 14353 7372 14358 7389
rect 14300 7355 14358 7372
rect 14300 7338 14336 7355
rect 14353 7338 14358 7355
rect 14300 7321 14358 7338
rect 14300 7304 14336 7321
rect 14353 7304 14358 7321
rect 14300 7287 14358 7304
rect 14300 7270 14336 7287
rect 14353 7270 14358 7287
rect 14300 7253 14358 7270
rect 14300 7236 14336 7253
rect 14353 7236 14358 7253
rect 14300 7219 14358 7236
rect 14300 7202 14336 7219
rect 14353 7202 14358 7219
rect 14300 7194 14358 7202
rect 14375 7389 14402 7412
rect 14986 7412 14990 7431
rect 15009 7412 15013 7431
rect 14375 7372 14380 7389
rect 14397 7372 14402 7389
rect 14375 7355 14402 7372
rect 14375 7338 14380 7355
rect 14397 7338 14402 7355
rect 14375 7321 14402 7338
rect 14375 7304 14380 7321
rect 14397 7304 14402 7321
rect 14375 7287 14402 7304
rect 14375 7270 14380 7287
rect 14397 7270 14402 7287
rect 14375 7253 14402 7270
rect 14375 7236 14380 7253
rect 14397 7236 14402 7253
rect 14375 7219 14402 7236
rect 14375 7202 14380 7219
rect 14397 7202 14402 7219
rect 14375 7194 14402 7202
rect 14419 7389 14477 7397
rect 14419 7372 14424 7389
rect 14441 7372 14477 7389
rect 14419 7355 14477 7372
rect 14419 7338 14424 7355
rect 14441 7338 14477 7355
rect 14419 7321 14477 7338
rect 14419 7304 14424 7321
rect 14441 7304 14477 7321
rect 14419 7287 14477 7304
rect 14419 7270 14424 7287
rect 14441 7270 14477 7287
rect 14419 7253 14477 7270
rect 14419 7236 14424 7253
rect 14441 7236 14477 7253
rect 14419 7219 14477 7236
rect 14419 7202 14424 7219
rect 14441 7202 14477 7219
rect 14419 7194 14477 7202
rect 14250 7117 14283 7125
rect 14250 7100 14258 7117
rect 14275 7100 14283 7117
rect 14250 7092 14283 7100
rect 14300 7107 14327 7194
rect 14349 7169 14382 7177
rect 14349 7152 14357 7169
rect 14374 7161 14382 7169
rect 14450 7161 14477 7194
rect 14374 7152 14477 7161
rect 14349 7144 14477 7152
rect 14395 7115 14428 7123
rect 14395 7107 14403 7115
rect 14300 7098 14403 7107
rect 14420 7098 14428 7115
rect 14300 7090 14428 7098
rect 13916 7079 13949 7087
rect 13916 7062 13924 7079
rect 13941 7062 13949 7079
rect 13916 7054 13949 7062
rect 14250 7063 14283 7071
rect 14250 7046 14258 7063
rect 14275 7046 14283 7063
rect 14250 7038 14283 7046
rect 14300 7021 14327 7090
rect 14450 7021 14477 7144
rect 14911 7389 14969 7397
rect 14911 7372 14947 7389
rect 14964 7372 14969 7389
rect 14911 7355 14969 7372
rect 14911 7338 14947 7355
rect 14964 7338 14969 7355
rect 14911 7321 14969 7338
rect 14911 7304 14947 7321
rect 14964 7304 14969 7321
rect 14911 7287 14969 7304
rect 14911 7270 14947 7287
rect 14964 7270 14969 7287
rect 14911 7253 14969 7270
rect 14911 7236 14947 7253
rect 14964 7236 14969 7253
rect 14911 7219 14969 7236
rect 14911 7202 14947 7219
rect 14964 7202 14969 7219
rect 14911 7194 14969 7202
rect 14986 7389 15013 7412
rect 15597 7412 15601 7431
rect 15620 7412 15624 7431
rect 14986 7372 14991 7389
rect 15008 7372 15013 7389
rect 14986 7355 15013 7372
rect 14986 7338 14991 7355
rect 15008 7338 15013 7355
rect 14986 7321 15013 7338
rect 14986 7304 14991 7321
rect 15008 7304 15013 7321
rect 14986 7287 15013 7304
rect 14986 7270 14991 7287
rect 15008 7270 15013 7287
rect 14986 7253 15013 7270
rect 14986 7236 14991 7253
rect 15008 7236 15013 7253
rect 14986 7219 15013 7236
rect 14986 7202 14991 7219
rect 15008 7202 15013 7219
rect 14986 7194 15013 7202
rect 15030 7389 15088 7397
rect 15030 7372 15035 7389
rect 15052 7372 15088 7389
rect 15030 7355 15088 7372
rect 15030 7338 15035 7355
rect 15052 7338 15088 7355
rect 15030 7321 15088 7338
rect 15030 7304 15035 7321
rect 15052 7304 15088 7321
rect 15030 7287 15088 7304
rect 15030 7270 15035 7287
rect 15052 7270 15088 7287
rect 15030 7253 15088 7270
rect 15030 7236 15035 7253
rect 15052 7236 15088 7253
rect 15030 7219 15088 7236
rect 15030 7202 15035 7219
rect 15052 7202 15088 7219
rect 15030 7194 15088 7202
rect 14861 7117 14894 7125
rect 14861 7100 14869 7117
rect 14886 7100 14894 7117
rect 14861 7092 14894 7100
rect 14911 7107 14938 7194
rect 14960 7169 14993 7177
rect 14960 7152 14968 7169
rect 14985 7161 14993 7169
rect 15061 7161 15088 7194
rect 14985 7152 15088 7161
rect 14960 7144 15088 7152
rect 15006 7115 15039 7123
rect 15006 7107 15014 7115
rect 14911 7098 15014 7107
rect 15031 7098 15039 7115
rect 14911 7090 15039 7098
rect 14494 7079 14527 7087
rect 14494 7062 14502 7079
rect 14519 7062 14527 7079
rect 14494 7054 14527 7062
rect 14861 7063 14894 7071
rect 14861 7046 14869 7063
rect 14886 7046 14894 7063
rect 14861 7038 14894 7046
rect 14911 7021 14938 7090
rect 15061 7021 15088 7144
rect 15522 7389 15580 7397
rect 15522 7372 15558 7389
rect 15575 7372 15580 7389
rect 15522 7355 15580 7372
rect 15522 7338 15558 7355
rect 15575 7338 15580 7355
rect 15522 7321 15580 7338
rect 15522 7304 15558 7321
rect 15575 7304 15580 7321
rect 15522 7287 15580 7304
rect 15522 7270 15558 7287
rect 15575 7270 15580 7287
rect 15522 7253 15580 7270
rect 15522 7236 15558 7253
rect 15575 7236 15580 7253
rect 15522 7219 15580 7236
rect 15522 7202 15558 7219
rect 15575 7202 15580 7219
rect 15522 7194 15580 7202
rect 15597 7389 15624 7412
rect 15597 7372 15602 7389
rect 15619 7372 15624 7389
rect 15597 7355 15624 7372
rect 15597 7338 15602 7355
rect 15619 7338 15624 7355
rect 15597 7321 15624 7338
rect 15597 7304 15602 7321
rect 15619 7304 15624 7321
rect 15597 7287 15624 7304
rect 15597 7270 15602 7287
rect 15619 7270 15624 7287
rect 15597 7253 15624 7270
rect 15597 7236 15602 7253
rect 15619 7236 15624 7253
rect 15597 7219 15624 7236
rect 15597 7202 15602 7219
rect 15619 7202 15624 7219
rect 15597 7194 15624 7202
rect 15641 7389 15699 7397
rect 15641 7372 15646 7389
rect 15663 7372 15699 7389
rect 15641 7355 15699 7372
rect 15641 7338 15646 7355
rect 15663 7338 15699 7355
rect 15641 7321 15699 7338
rect 15641 7304 15646 7321
rect 15663 7304 15699 7321
rect 15641 7287 15699 7304
rect 15641 7270 15646 7287
rect 15663 7270 15699 7287
rect 15641 7253 15699 7270
rect 15641 7236 15646 7253
rect 15663 7236 15699 7253
rect 15641 7219 15699 7236
rect 15641 7202 15646 7219
rect 15663 7202 15699 7219
rect 15641 7194 15699 7202
rect 15472 7117 15505 7125
rect 15472 7100 15480 7117
rect 15497 7100 15505 7117
rect 15472 7092 15505 7100
rect 15522 7107 15549 7194
rect 15571 7169 15604 7177
rect 15571 7152 15579 7169
rect 15596 7161 15604 7169
rect 15672 7161 15699 7194
rect 15596 7152 15699 7161
rect 15571 7144 15699 7152
rect 15617 7115 15650 7123
rect 15617 7107 15625 7115
rect 15522 7098 15625 7107
rect 15642 7098 15650 7115
rect 15522 7090 15650 7098
rect 15105 7079 15138 7087
rect 15105 7062 15113 7079
rect 15130 7062 15138 7079
rect 15105 7054 15138 7062
rect 15472 7063 15505 7071
rect 15472 7046 15480 7063
rect 15497 7046 15505 7063
rect 15472 7038 15505 7046
rect 15522 7021 15549 7090
rect 15672 7021 15699 7144
rect 15716 7079 15749 7087
rect 15716 7062 15724 7079
rect 15741 7062 15749 7079
rect 15716 7054 15749 7062
rect 12451 7013 12478 7021
rect 12451 6996 12456 7013
rect 12473 6996 12478 7013
rect 12451 6979 12478 6996
rect 12451 6962 12456 6979
rect 12473 6962 12478 6979
rect 12451 6945 12478 6962
rect 12451 6928 12456 6945
rect 12473 6928 12478 6945
rect 12451 6920 12478 6928
rect 12500 7013 12558 7021
rect 12500 6996 12536 7013
rect 12553 6996 12558 7013
rect 12500 6979 12558 6996
rect 12500 6962 12536 6979
rect 12553 6962 12558 6979
rect 12500 6945 12558 6962
rect 12500 6928 12536 6945
rect 12553 6928 12558 6945
rect 12500 6920 12558 6928
rect 12575 7013 12602 7021
rect 12575 6996 12580 7013
rect 12597 6996 12602 7013
rect 12575 6979 12602 6996
rect 12575 6962 12580 6979
rect 12597 6962 12602 6979
rect 12575 6945 12602 6962
rect 12575 6928 12580 6945
rect 12597 6928 12602 6945
rect 12575 6905 12602 6928
rect 12619 7013 12677 7021
rect 12619 6996 12624 7013
rect 12641 6996 12677 7013
rect 12619 6979 12677 6996
rect 12619 6962 12624 6979
rect 12641 6962 12677 6979
rect 12619 6945 12677 6962
rect 12619 6928 12624 6945
rect 12641 6928 12677 6945
rect 12619 6920 12677 6928
rect 12699 7013 12726 7021
rect 12699 6996 12704 7013
rect 12721 6996 12726 7013
rect 12699 6979 12726 6996
rect 12699 6962 12704 6979
rect 12721 6962 12726 6979
rect 12699 6945 12726 6962
rect 12699 6928 12704 6945
rect 12721 6928 12726 6945
rect 12699 6920 12726 6928
rect 13062 7013 13089 7021
rect 13062 6996 13067 7013
rect 13084 6996 13089 7013
rect 13062 6979 13089 6996
rect 13062 6962 13067 6979
rect 13084 6962 13089 6979
rect 13062 6945 13089 6962
rect 13062 6928 13067 6945
rect 13084 6928 13089 6945
rect 13062 6920 13089 6928
rect 13111 7013 13169 7021
rect 13111 6996 13147 7013
rect 13164 6996 13169 7013
rect 13111 6979 13169 6996
rect 13111 6962 13147 6979
rect 13164 6962 13169 6979
rect 13111 6945 13169 6962
rect 13111 6928 13147 6945
rect 13164 6928 13169 6945
rect 13111 6920 13169 6928
rect 13186 7013 13213 7021
rect 13186 6996 13191 7013
rect 13208 6996 13213 7013
rect 13186 6979 13213 6996
rect 13186 6962 13191 6979
rect 13208 6962 13213 6979
rect 13186 6945 13213 6962
rect 13186 6928 13191 6945
rect 13208 6928 13213 6945
rect 12575 6886 12579 6905
rect 12598 6886 12602 6905
rect 13186 6905 13213 6928
rect 13230 7013 13288 7021
rect 13230 6996 13235 7013
rect 13252 6996 13288 7013
rect 13230 6979 13288 6996
rect 13230 6962 13235 6979
rect 13252 6962 13288 6979
rect 13230 6945 13288 6962
rect 13230 6928 13235 6945
rect 13252 6928 13288 6945
rect 13230 6920 13288 6928
rect 13310 7013 13337 7021
rect 13310 6996 13315 7013
rect 13332 6996 13337 7013
rect 13310 6979 13337 6996
rect 13310 6962 13315 6979
rect 13332 6962 13337 6979
rect 13310 6945 13337 6962
rect 13310 6928 13315 6945
rect 13332 6928 13337 6945
rect 13310 6920 13337 6928
rect 13673 7013 13700 7021
rect 13673 6996 13678 7013
rect 13695 6996 13700 7013
rect 13673 6979 13700 6996
rect 13673 6962 13678 6979
rect 13695 6962 13700 6979
rect 13673 6945 13700 6962
rect 13673 6928 13678 6945
rect 13695 6928 13700 6945
rect 13673 6920 13700 6928
rect 13722 7013 13780 7021
rect 13722 6996 13758 7013
rect 13775 6996 13780 7013
rect 13722 6979 13780 6996
rect 13722 6962 13758 6979
rect 13775 6962 13780 6979
rect 13722 6945 13780 6962
rect 13722 6928 13758 6945
rect 13775 6928 13780 6945
rect 13722 6920 13780 6928
rect 13797 7013 13824 7021
rect 13797 6996 13802 7013
rect 13819 6996 13824 7013
rect 13797 6979 13824 6996
rect 13797 6962 13802 6979
rect 13819 6962 13824 6979
rect 13797 6945 13824 6962
rect 13797 6928 13802 6945
rect 13819 6928 13824 6945
rect 13186 6886 13190 6905
rect 13209 6886 13213 6905
rect 13797 6905 13824 6928
rect 13841 7013 13899 7021
rect 13841 6996 13846 7013
rect 13863 6996 13899 7013
rect 13841 6979 13899 6996
rect 13841 6962 13846 6979
rect 13863 6962 13899 6979
rect 13841 6945 13899 6962
rect 13841 6928 13846 6945
rect 13863 6928 13899 6945
rect 13841 6920 13899 6928
rect 13921 7013 13948 7021
rect 13921 6996 13926 7013
rect 13943 6996 13948 7013
rect 13921 6979 13948 6996
rect 13921 6962 13926 6979
rect 13943 6962 13948 6979
rect 13921 6945 13948 6962
rect 13921 6928 13926 6945
rect 13943 6928 13948 6945
rect 13921 6920 13948 6928
rect 14251 7013 14278 7021
rect 14251 6996 14256 7013
rect 14273 6996 14278 7013
rect 14251 6979 14278 6996
rect 14251 6962 14256 6979
rect 14273 6962 14278 6979
rect 14251 6945 14278 6962
rect 14251 6928 14256 6945
rect 14273 6928 14278 6945
rect 14251 6920 14278 6928
rect 14300 7013 14358 7021
rect 14300 6996 14336 7013
rect 14353 6996 14358 7013
rect 14300 6979 14358 6996
rect 14300 6962 14336 6979
rect 14353 6962 14358 6979
rect 14300 6945 14358 6962
rect 14300 6928 14336 6945
rect 14353 6928 14358 6945
rect 14300 6920 14358 6928
rect 14375 7013 14402 7021
rect 14375 6996 14380 7013
rect 14397 6996 14402 7013
rect 14375 6979 14402 6996
rect 14375 6962 14380 6979
rect 14397 6962 14402 6979
rect 14375 6945 14402 6962
rect 14375 6928 14380 6945
rect 14397 6928 14402 6945
rect 13797 6886 13801 6905
rect 13820 6886 13824 6905
rect 14375 6905 14402 6928
rect 14419 7013 14477 7021
rect 14419 6996 14424 7013
rect 14441 6996 14477 7013
rect 14419 6979 14477 6996
rect 14419 6962 14424 6979
rect 14441 6962 14477 6979
rect 14419 6945 14477 6962
rect 14419 6928 14424 6945
rect 14441 6928 14477 6945
rect 14419 6920 14477 6928
rect 14499 7013 14526 7021
rect 14499 6996 14504 7013
rect 14521 6996 14526 7013
rect 14499 6979 14526 6996
rect 14499 6962 14504 6979
rect 14521 6962 14526 6979
rect 14499 6945 14526 6962
rect 14499 6928 14504 6945
rect 14521 6928 14526 6945
rect 14499 6920 14526 6928
rect 14862 7013 14889 7021
rect 14862 6996 14867 7013
rect 14884 6996 14889 7013
rect 14862 6979 14889 6996
rect 14862 6962 14867 6979
rect 14884 6962 14889 6979
rect 14862 6945 14889 6962
rect 14862 6928 14867 6945
rect 14884 6928 14889 6945
rect 14862 6920 14889 6928
rect 14911 7013 14969 7021
rect 14911 6996 14947 7013
rect 14964 6996 14969 7013
rect 14911 6979 14969 6996
rect 14911 6962 14947 6979
rect 14964 6962 14969 6979
rect 14911 6945 14969 6962
rect 14911 6928 14947 6945
rect 14964 6928 14969 6945
rect 14911 6920 14969 6928
rect 14986 7013 15013 7021
rect 14986 6996 14991 7013
rect 15008 6996 15013 7013
rect 14986 6979 15013 6996
rect 14986 6962 14991 6979
rect 15008 6962 15013 6979
rect 14986 6945 15013 6962
rect 14986 6928 14991 6945
rect 15008 6928 15013 6945
rect 14375 6886 14379 6905
rect 14398 6886 14402 6905
rect 14986 6905 15013 6928
rect 15030 7013 15088 7021
rect 15030 6996 15035 7013
rect 15052 6996 15088 7013
rect 15030 6979 15088 6996
rect 15030 6962 15035 6979
rect 15052 6962 15088 6979
rect 15030 6945 15088 6962
rect 15030 6928 15035 6945
rect 15052 6928 15088 6945
rect 15030 6920 15088 6928
rect 15110 7013 15137 7021
rect 15110 6996 15115 7013
rect 15132 6996 15137 7013
rect 15110 6979 15137 6996
rect 15110 6962 15115 6979
rect 15132 6962 15137 6979
rect 15110 6945 15137 6962
rect 15110 6928 15115 6945
rect 15132 6928 15137 6945
rect 15110 6920 15137 6928
rect 15473 7013 15500 7021
rect 15473 6996 15478 7013
rect 15495 6996 15500 7013
rect 15473 6979 15500 6996
rect 15473 6962 15478 6979
rect 15495 6962 15500 6979
rect 15473 6945 15500 6962
rect 15473 6928 15478 6945
rect 15495 6928 15500 6945
rect 15473 6920 15500 6928
rect 15522 7013 15580 7021
rect 15522 6996 15558 7013
rect 15575 6996 15580 7013
rect 15522 6979 15580 6996
rect 15522 6962 15558 6979
rect 15575 6962 15580 6979
rect 15522 6945 15580 6962
rect 15522 6928 15558 6945
rect 15575 6928 15580 6945
rect 15522 6920 15580 6928
rect 15597 7013 15624 7021
rect 15597 6996 15602 7013
rect 15619 6996 15624 7013
rect 15597 6979 15624 6996
rect 15597 6962 15602 6979
rect 15619 6962 15624 6979
rect 15597 6945 15624 6962
rect 15597 6928 15602 6945
rect 15619 6928 15624 6945
rect 14986 6886 14990 6905
rect 15009 6886 15013 6905
rect 15597 6905 15624 6928
rect 15641 7013 15699 7021
rect 15641 6996 15646 7013
rect 15663 6996 15699 7013
rect 15641 6979 15699 6996
rect 15641 6962 15646 6979
rect 15663 6962 15699 6979
rect 15641 6945 15699 6962
rect 15641 6928 15646 6945
rect 15663 6928 15699 6945
rect 15641 6920 15699 6928
rect 15721 7013 15748 7021
rect 15721 6996 15726 7013
rect 15743 6996 15748 7013
rect 15721 6979 15748 6996
rect 15721 6962 15726 6979
rect 15743 6962 15748 6979
rect 15721 6945 15748 6962
rect 15721 6928 15726 6945
rect 15743 6928 15748 6945
rect 15721 6920 15748 6928
rect 15597 6886 15601 6905
rect 15620 6886 15624 6905
rect 12575 6772 12579 6791
rect 12598 6772 12602 6791
rect 12500 6749 12558 6757
rect 12500 6732 12536 6749
rect 12553 6732 12558 6749
rect 12500 6715 12558 6732
rect 12500 6698 12536 6715
rect 12553 6698 12558 6715
rect 12500 6681 12558 6698
rect 12500 6664 12536 6681
rect 12553 6664 12558 6681
rect 12500 6647 12558 6664
rect 12500 6630 12536 6647
rect 12553 6630 12558 6647
rect 12500 6613 12558 6630
rect 12500 6596 12536 6613
rect 12553 6596 12558 6613
rect 12500 6579 12558 6596
rect 12500 6562 12536 6579
rect 12553 6562 12558 6579
rect 12500 6554 12558 6562
rect 12575 6749 12602 6772
rect 13186 6772 13190 6791
rect 13209 6772 13213 6791
rect 12575 6732 12580 6749
rect 12597 6732 12602 6749
rect 12575 6715 12602 6732
rect 12575 6698 12580 6715
rect 12597 6698 12602 6715
rect 12575 6681 12602 6698
rect 12575 6664 12580 6681
rect 12597 6664 12602 6681
rect 12575 6647 12602 6664
rect 12575 6630 12580 6647
rect 12597 6630 12602 6647
rect 12575 6613 12602 6630
rect 12575 6596 12580 6613
rect 12597 6596 12602 6613
rect 12575 6579 12602 6596
rect 12575 6562 12580 6579
rect 12597 6562 12602 6579
rect 12575 6554 12602 6562
rect 12619 6749 12677 6757
rect 12619 6732 12624 6749
rect 12641 6732 12677 6749
rect 12619 6715 12677 6732
rect 12619 6698 12624 6715
rect 12641 6698 12677 6715
rect 12619 6681 12677 6698
rect 12619 6664 12624 6681
rect 12641 6664 12677 6681
rect 12619 6647 12677 6664
rect 12619 6630 12624 6647
rect 12641 6630 12677 6647
rect 12619 6613 12677 6630
rect 12619 6596 12624 6613
rect 12641 6596 12677 6613
rect 12619 6579 12677 6596
rect 12619 6562 12624 6579
rect 12641 6562 12677 6579
rect 12619 6554 12677 6562
rect 12450 6477 12483 6485
rect 12450 6460 12458 6477
rect 12475 6460 12483 6477
rect 12450 6452 12483 6460
rect 12500 6467 12527 6554
rect 12549 6529 12582 6537
rect 12549 6512 12557 6529
rect 12574 6521 12582 6529
rect 12650 6521 12677 6554
rect 12574 6512 12677 6521
rect 12549 6504 12677 6512
rect 12595 6475 12628 6483
rect 12595 6467 12603 6475
rect 12500 6458 12603 6467
rect 12620 6458 12628 6475
rect 12500 6450 12628 6458
rect 12450 6423 12483 6431
rect 12450 6406 12458 6423
rect 12475 6406 12483 6423
rect 12450 6398 12483 6406
rect 12500 6381 12527 6450
rect 12650 6381 12677 6504
rect 13111 6749 13169 6757
rect 13111 6732 13147 6749
rect 13164 6732 13169 6749
rect 13111 6715 13169 6732
rect 13111 6698 13147 6715
rect 13164 6698 13169 6715
rect 13111 6681 13169 6698
rect 13111 6664 13147 6681
rect 13164 6664 13169 6681
rect 13111 6647 13169 6664
rect 13111 6630 13147 6647
rect 13164 6630 13169 6647
rect 13111 6613 13169 6630
rect 13111 6596 13147 6613
rect 13164 6596 13169 6613
rect 13111 6579 13169 6596
rect 13111 6562 13147 6579
rect 13164 6562 13169 6579
rect 13111 6554 13169 6562
rect 13186 6749 13213 6772
rect 13797 6772 13801 6791
rect 13820 6772 13824 6791
rect 13186 6732 13191 6749
rect 13208 6732 13213 6749
rect 13186 6715 13213 6732
rect 13186 6698 13191 6715
rect 13208 6698 13213 6715
rect 13186 6681 13213 6698
rect 13186 6664 13191 6681
rect 13208 6664 13213 6681
rect 13186 6647 13213 6664
rect 13186 6630 13191 6647
rect 13208 6630 13213 6647
rect 13186 6613 13213 6630
rect 13186 6596 13191 6613
rect 13208 6596 13213 6613
rect 13186 6579 13213 6596
rect 13186 6562 13191 6579
rect 13208 6562 13213 6579
rect 13186 6554 13213 6562
rect 13230 6749 13288 6757
rect 13230 6732 13235 6749
rect 13252 6732 13288 6749
rect 13230 6715 13288 6732
rect 13230 6698 13235 6715
rect 13252 6698 13288 6715
rect 13230 6681 13288 6698
rect 13230 6664 13235 6681
rect 13252 6664 13288 6681
rect 13230 6647 13288 6664
rect 13230 6630 13235 6647
rect 13252 6630 13288 6647
rect 13230 6613 13288 6630
rect 13230 6596 13235 6613
rect 13252 6596 13288 6613
rect 13230 6579 13288 6596
rect 13230 6562 13235 6579
rect 13252 6562 13288 6579
rect 13230 6554 13288 6562
rect 13061 6477 13094 6485
rect 13061 6460 13069 6477
rect 13086 6460 13094 6477
rect 13061 6452 13094 6460
rect 13111 6467 13138 6554
rect 13160 6529 13193 6537
rect 13160 6512 13168 6529
rect 13185 6521 13193 6529
rect 13261 6521 13288 6554
rect 13185 6512 13288 6521
rect 13160 6504 13288 6512
rect 13206 6475 13239 6483
rect 13206 6467 13214 6475
rect 13111 6458 13214 6467
rect 13231 6458 13239 6475
rect 13111 6450 13239 6458
rect 12694 6439 12727 6447
rect 12694 6422 12702 6439
rect 12719 6422 12727 6439
rect 12694 6414 12727 6422
rect 13061 6423 13094 6431
rect 13061 6406 13069 6423
rect 13086 6406 13094 6423
rect 13061 6398 13094 6406
rect 13111 6381 13138 6450
rect 13261 6381 13288 6504
rect 13722 6749 13780 6757
rect 13722 6732 13758 6749
rect 13775 6732 13780 6749
rect 13722 6715 13780 6732
rect 13722 6698 13758 6715
rect 13775 6698 13780 6715
rect 13722 6681 13780 6698
rect 13722 6664 13758 6681
rect 13775 6664 13780 6681
rect 13722 6647 13780 6664
rect 13722 6630 13758 6647
rect 13775 6630 13780 6647
rect 13722 6613 13780 6630
rect 13722 6596 13758 6613
rect 13775 6596 13780 6613
rect 13722 6579 13780 6596
rect 13722 6562 13758 6579
rect 13775 6562 13780 6579
rect 13722 6554 13780 6562
rect 13797 6749 13824 6772
rect 14375 6772 14379 6791
rect 14398 6772 14402 6791
rect 13797 6732 13802 6749
rect 13819 6732 13824 6749
rect 13797 6715 13824 6732
rect 13797 6698 13802 6715
rect 13819 6698 13824 6715
rect 13797 6681 13824 6698
rect 13797 6664 13802 6681
rect 13819 6664 13824 6681
rect 13797 6647 13824 6664
rect 13797 6630 13802 6647
rect 13819 6630 13824 6647
rect 13797 6613 13824 6630
rect 13797 6596 13802 6613
rect 13819 6596 13824 6613
rect 13797 6579 13824 6596
rect 13797 6562 13802 6579
rect 13819 6562 13824 6579
rect 13797 6554 13824 6562
rect 13841 6749 13899 6757
rect 13841 6732 13846 6749
rect 13863 6732 13899 6749
rect 13841 6715 13899 6732
rect 13841 6698 13846 6715
rect 13863 6698 13899 6715
rect 13841 6681 13899 6698
rect 13841 6664 13846 6681
rect 13863 6664 13899 6681
rect 13841 6647 13899 6664
rect 13841 6630 13846 6647
rect 13863 6630 13899 6647
rect 13841 6613 13899 6630
rect 13841 6596 13846 6613
rect 13863 6596 13899 6613
rect 13841 6579 13899 6596
rect 13841 6562 13846 6579
rect 13863 6562 13899 6579
rect 13841 6554 13899 6562
rect 13672 6477 13705 6485
rect 13672 6460 13680 6477
rect 13697 6460 13705 6477
rect 13672 6452 13705 6460
rect 13722 6467 13749 6554
rect 13771 6529 13804 6537
rect 13771 6512 13779 6529
rect 13796 6521 13804 6529
rect 13872 6521 13899 6554
rect 13796 6512 13899 6521
rect 13771 6504 13899 6512
rect 13817 6475 13850 6483
rect 13817 6467 13825 6475
rect 13722 6458 13825 6467
rect 13842 6458 13850 6475
rect 13722 6450 13850 6458
rect 13305 6439 13338 6447
rect 13305 6422 13313 6439
rect 13330 6422 13338 6439
rect 13305 6414 13338 6422
rect 13672 6423 13705 6431
rect 13672 6406 13680 6423
rect 13697 6406 13705 6423
rect 13672 6398 13705 6406
rect 13722 6381 13749 6450
rect 13872 6381 13899 6504
rect 14300 6749 14358 6757
rect 14300 6732 14336 6749
rect 14353 6732 14358 6749
rect 14300 6715 14358 6732
rect 14300 6698 14336 6715
rect 14353 6698 14358 6715
rect 14300 6681 14358 6698
rect 14300 6664 14336 6681
rect 14353 6664 14358 6681
rect 14300 6647 14358 6664
rect 14300 6630 14336 6647
rect 14353 6630 14358 6647
rect 14300 6613 14358 6630
rect 14300 6596 14336 6613
rect 14353 6596 14358 6613
rect 14300 6579 14358 6596
rect 14300 6562 14336 6579
rect 14353 6562 14358 6579
rect 14300 6554 14358 6562
rect 14375 6749 14402 6772
rect 14986 6772 14990 6791
rect 15009 6772 15013 6791
rect 14375 6732 14380 6749
rect 14397 6732 14402 6749
rect 14375 6715 14402 6732
rect 14375 6698 14380 6715
rect 14397 6698 14402 6715
rect 14375 6681 14402 6698
rect 14375 6664 14380 6681
rect 14397 6664 14402 6681
rect 14375 6647 14402 6664
rect 14375 6630 14380 6647
rect 14397 6630 14402 6647
rect 14375 6613 14402 6630
rect 14375 6596 14380 6613
rect 14397 6596 14402 6613
rect 14375 6579 14402 6596
rect 14375 6562 14380 6579
rect 14397 6562 14402 6579
rect 14375 6554 14402 6562
rect 14419 6749 14477 6757
rect 14419 6732 14424 6749
rect 14441 6732 14477 6749
rect 14419 6715 14477 6732
rect 14419 6698 14424 6715
rect 14441 6698 14477 6715
rect 14419 6681 14477 6698
rect 14419 6664 14424 6681
rect 14441 6664 14477 6681
rect 14419 6647 14477 6664
rect 14419 6630 14424 6647
rect 14441 6630 14477 6647
rect 14419 6613 14477 6630
rect 14419 6596 14424 6613
rect 14441 6596 14477 6613
rect 14419 6579 14477 6596
rect 14419 6562 14424 6579
rect 14441 6562 14477 6579
rect 14419 6554 14477 6562
rect 14250 6477 14283 6485
rect 14250 6460 14258 6477
rect 14275 6460 14283 6477
rect 14250 6452 14283 6460
rect 14300 6467 14327 6554
rect 14349 6529 14382 6537
rect 14349 6512 14357 6529
rect 14374 6521 14382 6529
rect 14450 6521 14477 6554
rect 14374 6512 14477 6521
rect 14349 6504 14477 6512
rect 14395 6475 14428 6483
rect 14395 6467 14403 6475
rect 14300 6458 14403 6467
rect 14420 6458 14428 6475
rect 14300 6450 14428 6458
rect 13916 6439 13949 6447
rect 13916 6422 13924 6439
rect 13941 6422 13949 6439
rect 13916 6414 13949 6422
rect 14250 6423 14283 6431
rect 14250 6406 14258 6423
rect 14275 6406 14283 6423
rect 14250 6398 14283 6406
rect 14300 6381 14327 6450
rect 14450 6381 14477 6504
rect 14911 6749 14969 6757
rect 14911 6732 14947 6749
rect 14964 6732 14969 6749
rect 14911 6715 14969 6732
rect 14911 6698 14947 6715
rect 14964 6698 14969 6715
rect 14911 6681 14969 6698
rect 14911 6664 14947 6681
rect 14964 6664 14969 6681
rect 14911 6647 14969 6664
rect 14911 6630 14947 6647
rect 14964 6630 14969 6647
rect 14911 6613 14969 6630
rect 14911 6596 14947 6613
rect 14964 6596 14969 6613
rect 14911 6579 14969 6596
rect 14911 6562 14947 6579
rect 14964 6562 14969 6579
rect 14911 6554 14969 6562
rect 14986 6749 15013 6772
rect 15597 6772 15601 6791
rect 15620 6772 15624 6791
rect 14986 6732 14991 6749
rect 15008 6732 15013 6749
rect 14986 6715 15013 6732
rect 14986 6698 14991 6715
rect 15008 6698 15013 6715
rect 14986 6681 15013 6698
rect 14986 6664 14991 6681
rect 15008 6664 15013 6681
rect 14986 6647 15013 6664
rect 14986 6630 14991 6647
rect 15008 6630 15013 6647
rect 14986 6613 15013 6630
rect 14986 6596 14991 6613
rect 15008 6596 15013 6613
rect 14986 6579 15013 6596
rect 14986 6562 14991 6579
rect 15008 6562 15013 6579
rect 14986 6554 15013 6562
rect 15030 6749 15088 6757
rect 15030 6732 15035 6749
rect 15052 6732 15088 6749
rect 15030 6715 15088 6732
rect 15030 6698 15035 6715
rect 15052 6698 15088 6715
rect 15030 6681 15088 6698
rect 15030 6664 15035 6681
rect 15052 6664 15088 6681
rect 15030 6647 15088 6664
rect 15030 6630 15035 6647
rect 15052 6630 15088 6647
rect 15030 6613 15088 6630
rect 15030 6596 15035 6613
rect 15052 6596 15088 6613
rect 15030 6579 15088 6596
rect 15030 6562 15035 6579
rect 15052 6562 15088 6579
rect 15030 6554 15088 6562
rect 14861 6477 14894 6485
rect 14861 6460 14869 6477
rect 14886 6460 14894 6477
rect 14861 6452 14894 6460
rect 14911 6467 14938 6554
rect 14960 6529 14993 6537
rect 14960 6512 14968 6529
rect 14985 6521 14993 6529
rect 15061 6521 15088 6554
rect 14985 6512 15088 6521
rect 14960 6504 15088 6512
rect 15006 6475 15039 6483
rect 15006 6467 15014 6475
rect 14911 6458 15014 6467
rect 15031 6458 15039 6475
rect 14911 6450 15039 6458
rect 14494 6439 14527 6447
rect 14494 6422 14502 6439
rect 14519 6422 14527 6439
rect 14494 6414 14527 6422
rect 14861 6423 14894 6431
rect 14861 6406 14869 6423
rect 14886 6406 14894 6423
rect 14861 6398 14894 6406
rect 14911 6381 14938 6450
rect 15061 6381 15088 6504
rect 15522 6749 15580 6757
rect 15522 6732 15558 6749
rect 15575 6732 15580 6749
rect 15522 6715 15580 6732
rect 15522 6698 15558 6715
rect 15575 6698 15580 6715
rect 15522 6681 15580 6698
rect 15522 6664 15558 6681
rect 15575 6664 15580 6681
rect 15522 6647 15580 6664
rect 15522 6630 15558 6647
rect 15575 6630 15580 6647
rect 15522 6613 15580 6630
rect 15522 6596 15558 6613
rect 15575 6596 15580 6613
rect 15522 6579 15580 6596
rect 15522 6562 15558 6579
rect 15575 6562 15580 6579
rect 15522 6554 15580 6562
rect 15597 6749 15624 6772
rect 15597 6732 15602 6749
rect 15619 6732 15624 6749
rect 15597 6715 15624 6732
rect 15597 6698 15602 6715
rect 15619 6698 15624 6715
rect 15597 6681 15624 6698
rect 15597 6664 15602 6681
rect 15619 6664 15624 6681
rect 15597 6647 15624 6664
rect 15597 6630 15602 6647
rect 15619 6630 15624 6647
rect 15597 6613 15624 6630
rect 15597 6596 15602 6613
rect 15619 6596 15624 6613
rect 15597 6579 15624 6596
rect 15597 6562 15602 6579
rect 15619 6562 15624 6579
rect 15597 6554 15624 6562
rect 15641 6749 15699 6757
rect 15641 6732 15646 6749
rect 15663 6732 15699 6749
rect 15641 6715 15699 6732
rect 15641 6698 15646 6715
rect 15663 6698 15699 6715
rect 15641 6681 15699 6698
rect 15641 6664 15646 6681
rect 15663 6664 15699 6681
rect 15641 6647 15699 6664
rect 15641 6630 15646 6647
rect 15663 6630 15699 6647
rect 15641 6613 15699 6630
rect 15641 6596 15646 6613
rect 15663 6596 15699 6613
rect 15641 6579 15699 6596
rect 15641 6562 15646 6579
rect 15663 6562 15699 6579
rect 15641 6554 15699 6562
rect 15472 6477 15505 6485
rect 15472 6460 15480 6477
rect 15497 6460 15505 6477
rect 15472 6452 15505 6460
rect 15522 6467 15549 6554
rect 15571 6529 15604 6537
rect 15571 6512 15579 6529
rect 15596 6521 15604 6529
rect 15672 6521 15699 6554
rect 15596 6512 15699 6521
rect 15571 6504 15699 6512
rect 15617 6475 15650 6483
rect 15617 6467 15625 6475
rect 15522 6458 15625 6467
rect 15642 6458 15650 6475
rect 15522 6450 15650 6458
rect 15105 6439 15138 6447
rect 15105 6422 15113 6439
rect 15130 6422 15138 6439
rect 15105 6414 15138 6422
rect 15472 6423 15505 6431
rect 15472 6406 15480 6423
rect 15497 6406 15505 6423
rect 15472 6398 15505 6406
rect 15522 6381 15549 6450
rect 15672 6381 15699 6504
rect 15716 6439 15749 6447
rect 15716 6422 15724 6439
rect 15741 6422 15749 6439
rect 15716 6414 15749 6422
rect 12451 6373 12478 6381
rect 12451 6356 12456 6373
rect 12473 6356 12478 6373
rect 12451 6339 12478 6356
rect 12451 6322 12456 6339
rect 12473 6322 12478 6339
rect 12451 6305 12478 6322
rect 12451 6288 12456 6305
rect 12473 6288 12478 6305
rect 12451 6280 12478 6288
rect 12500 6373 12558 6381
rect 12500 6356 12536 6373
rect 12553 6356 12558 6373
rect 12500 6339 12558 6356
rect 12500 6322 12536 6339
rect 12553 6322 12558 6339
rect 12500 6305 12558 6322
rect 12500 6288 12536 6305
rect 12553 6288 12558 6305
rect 12500 6280 12558 6288
rect 12575 6373 12602 6381
rect 12575 6356 12580 6373
rect 12597 6356 12602 6373
rect 12575 6339 12602 6356
rect 12575 6322 12580 6339
rect 12597 6322 12602 6339
rect 12575 6305 12602 6322
rect 12575 6288 12580 6305
rect 12597 6288 12602 6305
rect 12575 6265 12602 6288
rect 12619 6373 12677 6381
rect 12619 6356 12624 6373
rect 12641 6356 12677 6373
rect 12619 6339 12677 6356
rect 12619 6322 12624 6339
rect 12641 6322 12677 6339
rect 12619 6305 12677 6322
rect 12619 6288 12624 6305
rect 12641 6288 12677 6305
rect 12619 6280 12677 6288
rect 12699 6373 12726 6381
rect 12699 6356 12704 6373
rect 12721 6356 12726 6373
rect 12699 6339 12726 6356
rect 12699 6322 12704 6339
rect 12721 6322 12726 6339
rect 12699 6305 12726 6322
rect 12699 6288 12704 6305
rect 12721 6288 12726 6305
rect 12699 6280 12726 6288
rect 13062 6373 13089 6381
rect 13062 6356 13067 6373
rect 13084 6356 13089 6373
rect 13062 6339 13089 6356
rect 13062 6322 13067 6339
rect 13084 6322 13089 6339
rect 13062 6305 13089 6322
rect 13062 6288 13067 6305
rect 13084 6288 13089 6305
rect 13062 6280 13089 6288
rect 13111 6373 13169 6381
rect 13111 6356 13147 6373
rect 13164 6356 13169 6373
rect 13111 6339 13169 6356
rect 13111 6322 13147 6339
rect 13164 6322 13169 6339
rect 13111 6305 13169 6322
rect 13111 6288 13147 6305
rect 13164 6288 13169 6305
rect 13111 6280 13169 6288
rect 13186 6373 13213 6381
rect 13186 6356 13191 6373
rect 13208 6356 13213 6373
rect 13186 6339 13213 6356
rect 13186 6322 13191 6339
rect 13208 6322 13213 6339
rect 13186 6305 13213 6322
rect 13186 6288 13191 6305
rect 13208 6288 13213 6305
rect 12575 6246 12579 6265
rect 12598 6246 12602 6265
rect 13186 6265 13213 6288
rect 13230 6373 13288 6381
rect 13230 6356 13235 6373
rect 13252 6356 13288 6373
rect 13230 6339 13288 6356
rect 13230 6322 13235 6339
rect 13252 6322 13288 6339
rect 13230 6305 13288 6322
rect 13230 6288 13235 6305
rect 13252 6288 13288 6305
rect 13230 6280 13288 6288
rect 13310 6373 13337 6381
rect 13310 6356 13315 6373
rect 13332 6356 13337 6373
rect 13310 6339 13337 6356
rect 13310 6322 13315 6339
rect 13332 6322 13337 6339
rect 13310 6305 13337 6322
rect 13310 6288 13315 6305
rect 13332 6288 13337 6305
rect 13310 6280 13337 6288
rect 13673 6373 13700 6381
rect 13673 6356 13678 6373
rect 13695 6356 13700 6373
rect 13673 6339 13700 6356
rect 13673 6322 13678 6339
rect 13695 6322 13700 6339
rect 13673 6305 13700 6322
rect 13673 6288 13678 6305
rect 13695 6288 13700 6305
rect 13673 6280 13700 6288
rect 13722 6373 13780 6381
rect 13722 6356 13758 6373
rect 13775 6356 13780 6373
rect 13722 6339 13780 6356
rect 13722 6322 13758 6339
rect 13775 6322 13780 6339
rect 13722 6305 13780 6322
rect 13722 6288 13758 6305
rect 13775 6288 13780 6305
rect 13722 6280 13780 6288
rect 13797 6373 13824 6381
rect 13797 6356 13802 6373
rect 13819 6356 13824 6373
rect 13797 6339 13824 6356
rect 13797 6322 13802 6339
rect 13819 6322 13824 6339
rect 13797 6305 13824 6322
rect 13797 6288 13802 6305
rect 13819 6288 13824 6305
rect 13186 6246 13190 6265
rect 13209 6246 13213 6265
rect 13797 6265 13824 6288
rect 13841 6373 13899 6381
rect 13841 6356 13846 6373
rect 13863 6356 13899 6373
rect 13841 6339 13899 6356
rect 13841 6322 13846 6339
rect 13863 6322 13899 6339
rect 13841 6305 13899 6322
rect 13841 6288 13846 6305
rect 13863 6288 13899 6305
rect 13841 6280 13899 6288
rect 13921 6373 13948 6381
rect 13921 6356 13926 6373
rect 13943 6356 13948 6373
rect 13921 6339 13948 6356
rect 13921 6322 13926 6339
rect 13943 6322 13948 6339
rect 13921 6305 13948 6322
rect 13921 6288 13926 6305
rect 13943 6288 13948 6305
rect 13921 6280 13948 6288
rect 14251 6373 14278 6381
rect 14251 6356 14256 6373
rect 14273 6356 14278 6373
rect 14251 6339 14278 6356
rect 14251 6322 14256 6339
rect 14273 6322 14278 6339
rect 14251 6305 14278 6322
rect 14251 6288 14256 6305
rect 14273 6288 14278 6305
rect 14251 6280 14278 6288
rect 14300 6373 14358 6381
rect 14300 6356 14336 6373
rect 14353 6356 14358 6373
rect 14300 6339 14358 6356
rect 14300 6322 14336 6339
rect 14353 6322 14358 6339
rect 14300 6305 14358 6322
rect 14300 6288 14336 6305
rect 14353 6288 14358 6305
rect 14300 6280 14358 6288
rect 14375 6373 14402 6381
rect 14375 6356 14380 6373
rect 14397 6356 14402 6373
rect 14375 6339 14402 6356
rect 14375 6322 14380 6339
rect 14397 6322 14402 6339
rect 14375 6305 14402 6322
rect 14375 6288 14380 6305
rect 14397 6288 14402 6305
rect 13797 6246 13801 6265
rect 13820 6246 13824 6265
rect 14375 6265 14402 6288
rect 14419 6373 14477 6381
rect 14419 6356 14424 6373
rect 14441 6356 14477 6373
rect 14419 6339 14477 6356
rect 14419 6322 14424 6339
rect 14441 6322 14477 6339
rect 14419 6305 14477 6322
rect 14419 6288 14424 6305
rect 14441 6288 14477 6305
rect 14419 6280 14477 6288
rect 14499 6373 14526 6381
rect 14499 6356 14504 6373
rect 14521 6356 14526 6373
rect 14499 6339 14526 6356
rect 14499 6322 14504 6339
rect 14521 6322 14526 6339
rect 14499 6305 14526 6322
rect 14499 6288 14504 6305
rect 14521 6288 14526 6305
rect 14499 6280 14526 6288
rect 14862 6373 14889 6381
rect 14862 6356 14867 6373
rect 14884 6356 14889 6373
rect 14862 6339 14889 6356
rect 14862 6322 14867 6339
rect 14884 6322 14889 6339
rect 14862 6305 14889 6322
rect 14862 6288 14867 6305
rect 14884 6288 14889 6305
rect 14862 6280 14889 6288
rect 14911 6373 14969 6381
rect 14911 6356 14947 6373
rect 14964 6356 14969 6373
rect 14911 6339 14969 6356
rect 14911 6322 14947 6339
rect 14964 6322 14969 6339
rect 14911 6305 14969 6322
rect 14911 6288 14947 6305
rect 14964 6288 14969 6305
rect 14911 6280 14969 6288
rect 14986 6373 15013 6381
rect 14986 6356 14991 6373
rect 15008 6356 15013 6373
rect 14986 6339 15013 6356
rect 14986 6322 14991 6339
rect 15008 6322 15013 6339
rect 14986 6305 15013 6322
rect 14986 6288 14991 6305
rect 15008 6288 15013 6305
rect 14375 6246 14379 6265
rect 14398 6246 14402 6265
rect 14986 6265 15013 6288
rect 15030 6373 15088 6381
rect 15030 6356 15035 6373
rect 15052 6356 15088 6373
rect 15030 6339 15088 6356
rect 15030 6322 15035 6339
rect 15052 6322 15088 6339
rect 15030 6305 15088 6322
rect 15030 6288 15035 6305
rect 15052 6288 15088 6305
rect 15030 6280 15088 6288
rect 15110 6373 15137 6381
rect 15110 6356 15115 6373
rect 15132 6356 15137 6373
rect 15110 6339 15137 6356
rect 15110 6322 15115 6339
rect 15132 6322 15137 6339
rect 15110 6305 15137 6322
rect 15110 6288 15115 6305
rect 15132 6288 15137 6305
rect 15110 6280 15137 6288
rect 15473 6373 15500 6381
rect 15473 6356 15478 6373
rect 15495 6356 15500 6373
rect 15473 6339 15500 6356
rect 15473 6322 15478 6339
rect 15495 6322 15500 6339
rect 15473 6305 15500 6322
rect 15473 6288 15478 6305
rect 15495 6288 15500 6305
rect 15473 6280 15500 6288
rect 15522 6373 15580 6381
rect 15522 6356 15558 6373
rect 15575 6356 15580 6373
rect 15522 6339 15580 6356
rect 15522 6322 15558 6339
rect 15575 6322 15580 6339
rect 15522 6305 15580 6322
rect 15522 6288 15558 6305
rect 15575 6288 15580 6305
rect 15522 6280 15580 6288
rect 15597 6373 15624 6381
rect 15597 6356 15602 6373
rect 15619 6356 15624 6373
rect 15597 6339 15624 6356
rect 15597 6322 15602 6339
rect 15619 6322 15624 6339
rect 15597 6305 15624 6322
rect 15597 6288 15602 6305
rect 15619 6288 15624 6305
rect 14986 6246 14990 6265
rect 15009 6246 15013 6265
rect 15597 6265 15624 6288
rect 15641 6373 15699 6381
rect 15641 6356 15646 6373
rect 15663 6356 15699 6373
rect 15641 6339 15699 6356
rect 15641 6322 15646 6339
rect 15663 6322 15699 6339
rect 15641 6305 15699 6322
rect 15641 6288 15646 6305
rect 15663 6288 15699 6305
rect 15641 6280 15699 6288
rect 15721 6373 15748 6381
rect 15721 6356 15726 6373
rect 15743 6356 15748 6373
rect 15721 6339 15748 6356
rect 15721 6322 15726 6339
rect 15743 6322 15748 6339
rect 15721 6305 15748 6322
rect 15721 6288 15726 6305
rect 15743 6288 15748 6305
rect 15721 6280 15748 6288
rect 15597 6246 15601 6265
rect 15620 6246 15624 6265
rect 12575 6122 12579 6141
rect 12598 6122 12602 6141
rect 12500 6099 12558 6107
rect 12500 6082 12536 6099
rect 12553 6082 12558 6099
rect 12500 6065 12558 6082
rect 12500 6048 12536 6065
rect 12553 6048 12558 6065
rect 12500 6031 12558 6048
rect 12500 6014 12536 6031
rect 12553 6014 12558 6031
rect 12500 5997 12558 6014
rect 12500 5980 12536 5997
rect 12553 5980 12558 5997
rect 12500 5963 12558 5980
rect 12500 5946 12536 5963
rect 12553 5946 12558 5963
rect 12500 5929 12558 5946
rect 12500 5912 12536 5929
rect 12553 5912 12558 5929
rect 12500 5904 12558 5912
rect 12575 6099 12602 6122
rect 13186 6122 13190 6141
rect 13209 6122 13213 6141
rect 12575 6082 12580 6099
rect 12597 6082 12602 6099
rect 12575 6065 12602 6082
rect 12575 6048 12580 6065
rect 12597 6048 12602 6065
rect 12575 6031 12602 6048
rect 12575 6014 12580 6031
rect 12597 6014 12602 6031
rect 12575 5997 12602 6014
rect 12575 5980 12580 5997
rect 12597 5980 12602 5997
rect 12575 5963 12602 5980
rect 12575 5946 12580 5963
rect 12597 5946 12602 5963
rect 12575 5929 12602 5946
rect 12575 5912 12580 5929
rect 12597 5912 12602 5929
rect 12575 5904 12602 5912
rect 12619 6099 12677 6107
rect 12619 6082 12624 6099
rect 12641 6082 12677 6099
rect 12619 6065 12677 6082
rect 12619 6048 12624 6065
rect 12641 6048 12677 6065
rect 12619 6031 12677 6048
rect 12619 6014 12624 6031
rect 12641 6014 12677 6031
rect 12619 5997 12677 6014
rect 12619 5980 12624 5997
rect 12641 5980 12677 5997
rect 12619 5963 12677 5980
rect 12619 5946 12624 5963
rect 12641 5946 12677 5963
rect 12619 5929 12677 5946
rect 12619 5912 12624 5929
rect 12641 5912 12677 5929
rect 12619 5904 12677 5912
rect 12450 5827 12483 5835
rect 12450 5810 12458 5827
rect 12475 5810 12483 5827
rect 12450 5802 12483 5810
rect 12500 5817 12527 5904
rect 12549 5879 12582 5887
rect 12549 5862 12557 5879
rect 12574 5871 12582 5879
rect 12650 5871 12677 5904
rect 12574 5862 12677 5871
rect 12549 5854 12677 5862
rect 12595 5825 12628 5833
rect 12595 5817 12603 5825
rect 12500 5808 12603 5817
rect 12620 5808 12628 5825
rect 12500 5800 12628 5808
rect 12450 5773 12483 5781
rect 12450 5756 12458 5773
rect 12475 5756 12483 5773
rect 12450 5748 12483 5756
rect 12500 5731 12527 5800
rect 12650 5731 12677 5854
rect 13111 6099 13169 6107
rect 13111 6082 13147 6099
rect 13164 6082 13169 6099
rect 13111 6065 13169 6082
rect 13111 6048 13147 6065
rect 13164 6048 13169 6065
rect 13111 6031 13169 6048
rect 13111 6014 13147 6031
rect 13164 6014 13169 6031
rect 13111 5997 13169 6014
rect 13111 5980 13147 5997
rect 13164 5980 13169 5997
rect 13111 5963 13169 5980
rect 13111 5946 13147 5963
rect 13164 5946 13169 5963
rect 13111 5929 13169 5946
rect 13111 5912 13147 5929
rect 13164 5912 13169 5929
rect 13111 5904 13169 5912
rect 13186 6099 13213 6122
rect 13797 6122 13801 6141
rect 13820 6122 13824 6141
rect 13186 6082 13191 6099
rect 13208 6082 13213 6099
rect 13186 6065 13213 6082
rect 13186 6048 13191 6065
rect 13208 6048 13213 6065
rect 13186 6031 13213 6048
rect 13186 6014 13191 6031
rect 13208 6014 13213 6031
rect 13186 5997 13213 6014
rect 13186 5980 13191 5997
rect 13208 5980 13213 5997
rect 13186 5963 13213 5980
rect 13186 5946 13191 5963
rect 13208 5946 13213 5963
rect 13186 5929 13213 5946
rect 13186 5912 13191 5929
rect 13208 5912 13213 5929
rect 13186 5904 13213 5912
rect 13230 6099 13288 6107
rect 13230 6082 13235 6099
rect 13252 6082 13288 6099
rect 13230 6065 13288 6082
rect 13230 6048 13235 6065
rect 13252 6048 13288 6065
rect 13230 6031 13288 6048
rect 13230 6014 13235 6031
rect 13252 6014 13288 6031
rect 13230 5997 13288 6014
rect 13230 5980 13235 5997
rect 13252 5980 13288 5997
rect 13230 5963 13288 5980
rect 13230 5946 13235 5963
rect 13252 5946 13288 5963
rect 13230 5929 13288 5946
rect 13230 5912 13235 5929
rect 13252 5912 13288 5929
rect 13230 5904 13288 5912
rect 13061 5827 13094 5835
rect 13061 5810 13069 5827
rect 13086 5810 13094 5827
rect 13061 5802 13094 5810
rect 13111 5817 13138 5904
rect 13160 5879 13193 5887
rect 13160 5862 13168 5879
rect 13185 5871 13193 5879
rect 13261 5871 13288 5904
rect 13185 5862 13288 5871
rect 13160 5854 13288 5862
rect 13206 5825 13239 5833
rect 13206 5817 13214 5825
rect 13111 5808 13214 5817
rect 13231 5808 13239 5825
rect 13111 5800 13239 5808
rect 12694 5789 12727 5797
rect 12694 5772 12702 5789
rect 12719 5772 12727 5789
rect 12694 5764 12727 5772
rect 13061 5773 13094 5781
rect 13061 5756 13069 5773
rect 13086 5756 13094 5773
rect 13061 5748 13094 5756
rect 13111 5731 13138 5800
rect 13261 5731 13288 5854
rect 13722 6099 13780 6107
rect 13722 6082 13758 6099
rect 13775 6082 13780 6099
rect 13722 6065 13780 6082
rect 13722 6048 13758 6065
rect 13775 6048 13780 6065
rect 13722 6031 13780 6048
rect 13722 6014 13758 6031
rect 13775 6014 13780 6031
rect 13722 5997 13780 6014
rect 13722 5980 13758 5997
rect 13775 5980 13780 5997
rect 13722 5963 13780 5980
rect 13722 5946 13758 5963
rect 13775 5946 13780 5963
rect 13722 5929 13780 5946
rect 13722 5912 13758 5929
rect 13775 5912 13780 5929
rect 13722 5904 13780 5912
rect 13797 6099 13824 6122
rect 14375 6122 14379 6141
rect 14398 6122 14402 6141
rect 13797 6082 13802 6099
rect 13819 6082 13824 6099
rect 13797 6065 13824 6082
rect 13797 6048 13802 6065
rect 13819 6048 13824 6065
rect 13797 6031 13824 6048
rect 13797 6014 13802 6031
rect 13819 6014 13824 6031
rect 13797 5997 13824 6014
rect 13797 5980 13802 5997
rect 13819 5980 13824 5997
rect 13797 5963 13824 5980
rect 13797 5946 13802 5963
rect 13819 5946 13824 5963
rect 13797 5929 13824 5946
rect 13797 5912 13802 5929
rect 13819 5912 13824 5929
rect 13797 5904 13824 5912
rect 13841 6099 13899 6107
rect 13841 6082 13846 6099
rect 13863 6082 13899 6099
rect 13841 6065 13899 6082
rect 13841 6048 13846 6065
rect 13863 6048 13899 6065
rect 13841 6031 13899 6048
rect 13841 6014 13846 6031
rect 13863 6014 13899 6031
rect 13841 5997 13899 6014
rect 13841 5980 13846 5997
rect 13863 5980 13899 5997
rect 13841 5963 13899 5980
rect 13841 5946 13846 5963
rect 13863 5946 13899 5963
rect 13841 5929 13899 5946
rect 13841 5912 13846 5929
rect 13863 5912 13899 5929
rect 13841 5904 13899 5912
rect 13672 5827 13705 5835
rect 13672 5810 13680 5827
rect 13697 5810 13705 5827
rect 13672 5802 13705 5810
rect 13722 5817 13749 5904
rect 13771 5879 13804 5887
rect 13771 5862 13779 5879
rect 13796 5871 13804 5879
rect 13872 5871 13899 5904
rect 13796 5862 13899 5871
rect 13771 5854 13899 5862
rect 13817 5825 13850 5833
rect 13817 5817 13825 5825
rect 13722 5808 13825 5817
rect 13842 5808 13850 5825
rect 13722 5800 13850 5808
rect 13305 5789 13338 5797
rect 13305 5772 13313 5789
rect 13330 5772 13338 5789
rect 13305 5764 13338 5772
rect 13672 5773 13705 5781
rect 13672 5756 13680 5773
rect 13697 5756 13705 5773
rect 13672 5748 13705 5756
rect 13722 5731 13749 5800
rect 13872 5731 13899 5854
rect 14300 6099 14358 6107
rect 14300 6082 14336 6099
rect 14353 6082 14358 6099
rect 14300 6065 14358 6082
rect 14300 6048 14336 6065
rect 14353 6048 14358 6065
rect 14300 6031 14358 6048
rect 14300 6014 14336 6031
rect 14353 6014 14358 6031
rect 14300 5997 14358 6014
rect 14300 5980 14336 5997
rect 14353 5980 14358 5997
rect 14300 5963 14358 5980
rect 14300 5946 14336 5963
rect 14353 5946 14358 5963
rect 14300 5929 14358 5946
rect 14300 5912 14336 5929
rect 14353 5912 14358 5929
rect 14300 5904 14358 5912
rect 14375 6099 14402 6122
rect 14986 6122 14990 6141
rect 15009 6122 15013 6141
rect 14375 6082 14380 6099
rect 14397 6082 14402 6099
rect 14375 6065 14402 6082
rect 14375 6048 14380 6065
rect 14397 6048 14402 6065
rect 14375 6031 14402 6048
rect 14375 6014 14380 6031
rect 14397 6014 14402 6031
rect 14375 5997 14402 6014
rect 14375 5980 14380 5997
rect 14397 5980 14402 5997
rect 14375 5963 14402 5980
rect 14375 5946 14380 5963
rect 14397 5946 14402 5963
rect 14375 5929 14402 5946
rect 14375 5912 14380 5929
rect 14397 5912 14402 5929
rect 14375 5904 14402 5912
rect 14419 6099 14477 6107
rect 14419 6082 14424 6099
rect 14441 6082 14477 6099
rect 14419 6065 14477 6082
rect 14419 6048 14424 6065
rect 14441 6048 14477 6065
rect 14419 6031 14477 6048
rect 14419 6014 14424 6031
rect 14441 6014 14477 6031
rect 14419 5997 14477 6014
rect 14419 5980 14424 5997
rect 14441 5980 14477 5997
rect 14419 5963 14477 5980
rect 14419 5946 14424 5963
rect 14441 5946 14477 5963
rect 14419 5929 14477 5946
rect 14419 5912 14424 5929
rect 14441 5912 14477 5929
rect 14419 5904 14477 5912
rect 14250 5827 14283 5835
rect 14250 5810 14258 5827
rect 14275 5810 14283 5827
rect 14250 5802 14283 5810
rect 14300 5817 14327 5904
rect 14349 5879 14382 5887
rect 14349 5862 14357 5879
rect 14374 5871 14382 5879
rect 14450 5871 14477 5904
rect 14374 5862 14477 5871
rect 14349 5854 14477 5862
rect 14395 5825 14428 5833
rect 14395 5817 14403 5825
rect 14300 5808 14403 5817
rect 14420 5808 14428 5825
rect 14300 5800 14428 5808
rect 13916 5789 13949 5797
rect 13916 5772 13924 5789
rect 13941 5772 13949 5789
rect 13916 5764 13949 5772
rect 14250 5773 14283 5781
rect 14250 5756 14258 5773
rect 14275 5756 14283 5773
rect 14250 5748 14283 5756
rect 14300 5731 14327 5800
rect 14450 5731 14477 5854
rect 14911 6099 14969 6107
rect 14911 6082 14947 6099
rect 14964 6082 14969 6099
rect 14911 6065 14969 6082
rect 14911 6048 14947 6065
rect 14964 6048 14969 6065
rect 14911 6031 14969 6048
rect 14911 6014 14947 6031
rect 14964 6014 14969 6031
rect 14911 5997 14969 6014
rect 14911 5980 14947 5997
rect 14964 5980 14969 5997
rect 14911 5963 14969 5980
rect 14911 5946 14947 5963
rect 14964 5946 14969 5963
rect 14911 5929 14969 5946
rect 14911 5912 14947 5929
rect 14964 5912 14969 5929
rect 14911 5904 14969 5912
rect 14986 6099 15013 6122
rect 15597 6122 15601 6141
rect 15620 6122 15624 6141
rect 14986 6082 14991 6099
rect 15008 6082 15013 6099
rect 14986 6065 15013 6082
rect 14986 6048 14991 6065
rect 15008 6048 15013 6065
rect 14986 6031 15013 6048
rect 14986 6014 14991 6031
rect 15008 6014 15013 6031
rect 14986 5997 15013 6014
rect 14986 5980 14991 5997
rect 15008 5980 15013 5997
rect 14986 5963 15013 5980
rect 14986 5946 14991 5963
rect 15008 5946 15013 5963
rect 14986 5929 15013 5946
rect 14986 5912 14991 5929
rect 15008 5912 15013 5929
rect 14986 5904 15013 5912
rect 15030 6099 15088 6107
rect 15030 6082 15035 6099
rect 15052 6082 15088 6099
rect 15030 6065 15088 6082
rect 15030 6048 15035 6065
rect 15052 6048 15088 6065
rect 15030 6031 15088 6048
rect 15030 6014 15035 6031
rect 15052 6014 15088 6031
rect 15030 5997 15088 6014
rect 15030 5980 15035 5997
rect 15052 5980 15088 5997
rect 15030 5963 15088 5980
rect 15030 5946 15035 5963
rect 15052 5946 15088 5963
rect 15030 5929 15088 5946
rect 15030 5912 15035 5929
rect 15052 5912 15088 5929
rect 15030 5904 15088 5912
rect 14861 5827 14894 5835
rect 14861 5810 14869 5827
rect 14886 5810 14894 5827
rect 14861 5802 14894 5810
rect 14911 5817 14938 5904
rect 14960 5879 14993 5887
rect 14960 5862 14968 5879
rect 14985 5871 14993 5879
rect 15061 5871 15088 5904
rect 14985 5862 15088 5871
rect 14960 5854 15088 5862
rect 15006 5825 15039 5833
rect 15006 5817 15014 5825
rect 14911 5808 15014 5817
rect 15031 5808 15039 5825
rect 14911 5800 15039 5808
rect 14494 5789 14527 5797
rect 14494 5772 14502 5789
rect 14519 5772 14527 5789
rect 14494 5764 14527 5772
rect 14861 5773 14894 5781
rect 14861 5756 14869 5773
rect 14886 5756 14894 5773
rect 14861 5748 14894 5756
rect 14911 5731 14938 5800
rect 15061 5731 15088 5854
rect 15522 6099 15580 6107
rect 15522 6082 15558 6099
rect 15575 6082 15580 6099
rect 15522 6065 15580 6082
rect 15522 6048 15558 6065
rect 15575 6048 15580 6065
rect 15522 6031 15580 6048
rect 15522 6014 15558 6031
rect 15575 6014 15580 6031
rect 15522 5997 15580 6014
rect 15522 5980 15558 5997
rect 15575 5980 15580 5997
rect 15522 5963 15580 5980
rect 15522 5946 15558 5963
rect 15575 5946 15580 5963
rect 15522 5929 15580 5946
rect 15522 5912 15558 5929
rect 15575 5912 15580 5929
rect 15522 5904 15580 5912
rect 15597 6099 15624 6122
rect 15597 6082 15602 6099
rect 15619 6082 15624 6099
rect 15597 6065 15624 6082
rect 15597 6048 15602 6065
rect 15619 6048 15624 6065
rect 15597 6031 15624 6048
rect 15597 6014 15602 6031
rect 15619 6014 15624 6031
rect 15597 5997 15624 6014
rect 15597 5980 15602 5997
rect 15619 5980 15624 5997
rect 15597 5963 15624 5980
rect 15597 5946 15602 5963
rect 15619 5946 15624 5963
rect 15597 5929 15624 5946
rect 15597 5912 15602 5929
rect 15619 5912 15624 5929
rect 15597 5904 15624 5912
rect 15641 6099 15699 6107
rect 15641 6082 15646 6099
rect 15663 6082 15699 6099
rect 15641 6065 15699 6082
rect 15641 6048 15646 6065
rect 15663 6048 15699 6065
rect 15641 6031 15699 6048
rect 15641 6014 15646 6031
rect 15663 6014 15699 6031
rect 15641 5997 15699 6014
rect 15641 5980 15646 5997
rect 15663 5980 15699 5997
rect 15641 5963 15699 5980
rect 15641 5946 15646 5963
rect 15663 5946 15699 5963
rect 15641 5929 15699 5946
rect 15641 5912 15646 5929
rect 15663 5912 15699 5929
rect 15641 5904 15699 5912
rect 15472 5827 15505 5835
rect 15472 5810 15480 5827
rect 15497 5810 15505 5827
rect 15472 5802 15505 5810
rect 15522 5817 15549 5904
rect 15571 5879 15604 5887
rect 15571 5862 15579 5879
rect 15596 5871 15604 5879
rect 15672 5871 15699 5904
rect 15596 5862 15699 5871
rect 15571 5854 15699 5862
rect 15617 5825 15650 5833
rect 15617 5817 15625 5825
rect 15522 5808 15625 5817
rect 15642 5808 15650 5825
rect 15522 5800 15650 5808
rect 15105 5789 15138 5797
rect 15105 5772 15113 5789
rect 15130 5772 15138 5789
rect 15105 5764 15138 5772
rect 15472 5773 15505 5781
rect 15472 5756 15480 5773
rect 15497 5756 15505 5773
rect 15472 5748 15505 5756
rect 15522 5731 15549 5800
rect 15672 5731 15699 5854
rect 15716 5789 15749 5797
rect 15716 5772 15724 5789
rect 15741 5772 15749 5789
rect 15716 5764 15749 5772
rect 12451 5723 12478 5731
rect 12451 5706 12456 5723
rect 12473 5706 12478 5723
rect 12451 5689 12478 5706
rect 12451 5672 12456 5689
rect 12473 5672 12478 5689
rect 12451 5655 12478 5672
rect 12451 5638 12456 5655
rect 12473 5638 12478 5655
rect 12451 5630 12478 5638
rect 12500 5723 12558 5731
rect 12500 5706 12536 5723
rect 12553 5706 12558 5723
rect 12500 5689 12558 5706
rect 12500 5672 12536 5689
rect 12553 5672 12558 5689
rect 12500 5655 12558 5672
rect 12500 5638 12536 5655
rect 12553 5638 12558 5655
rect 12500 5630 12558 5638
rect 12575 5723 12602 5731
rect 12575 5706 12580 5723
rect 12597 5706 12602 5723
rect 12575 5689 12602 5706
rect 12575 5672 12580 5689
rect 12597 5672 12602 5689
rect 12575 5655 12602 5672
rect 12575 5638 12580 5655
rect 12597 5638 12602 5655
rect 12575 5615 12602 5638
rect 12619 5723 12677 5731
rect 12619 5706 12624 5723
rect 12641 5706 12677 5723
rect 12619 5689 12677 5706
rect 12619 5672 12624 5689
rect 12641 5672 12677 5689
rect 12619 5655 12677 5672
rect 12619 5638 12624 5655
rect 12641 5638 12677 5655
rect 12619 5630 12677 5638
rect 12699 5723 12726 5731
rect 12699 5706 12704 5723
rect 12721 5706 12726 5723
rect 12699 5689 12726 5706
rect 12699 5672 12704 5689
rect 12721 5672 12726 5689
rect 12699 5655 12726 5672
rect 12699 5638 12704 5655
rect 12721 5638 12726 5655
rect 12699 5630 12726 5638
rect 13062 5723 13089 5731
rect 13062 5706 13067 5723
rect 13084 5706 13089 5723
rect 13062 5689 13089 5706
rect 13062 5672 13067 5689
rect 13084 5672 13089 5689
rect 13062 5655 13089 5672
rect 13062 5638 13067 5655
rect 13084 5638 13089 5655
rect 13062 5630 13089 5638
rect 13111 5723 13169 5731
rect 13111 5706 13147 5723
rect 13164 5706 13169 5723
rect 13111 5689 13169 5706
rect 13111 5672 13147 5689
rect 13164 5672 13169 5689
rect 13111 5655 13169 5672
rect 13111 5638 13147 5655
rect 13164 5638 13169 5655
rect 13111 5630 13169 5638
rect 13186 5723 13213 5731
rect 13186 5706 13191 5723
rect 13208 5706 13213 5723
rect 13186 5689 13213 5706
rect 13186 5672 13191 5689
rect 13208 5672 13213 5689
rect 13186 5655 13213 5672
rect 13186 5638 13191 5655
rect 13208 5638 13213 5655
rect 12575 5596 12579 5615
rect 12598 5596 12602 5615
rect 13186 5615 13213 5638
rect 13230 5723 13288 5731
rect 13230 5706 13235 5723
rect 13252 5706 13288 5723
rect 13230 5689 13288 5706
rect 13230 5672 13235 5689
rect 13252 5672 13288 5689
rect 13230 5655 13288 5672
rect 13230 5638 13235 5655
rect 13252 5638 13288 5655
rect 13230 5630 13288 5638
rect 13310 5723 13337 5731
rect 13310 5706 13315 5723
rect 13332 5706 13337 5723
rect 13310 5689 13337 5706
rect 13310 5672 13315 5689
rect 13332 5672 13337 5689
rect 13310 5655 13337 5672
rect 13310 5638 13315 5655
rect 13332 5638 13337 5655
rect 13310 5630 13337 5638
rect 13673 5723 13700 5731
rect 13673 5706 13678 5723
rect 13695 5706 13700 5723
rect 13673 5689 13700 5706
rect 13673 5672 13678 5689
rect 13695 5672 13700 5689
rect 13673 5655 13700 5672
rect 13673 5638 13678 5655
rect 13695 5638 13700 5655
rect 13673 5630 13700 5638
rect 13722 5723 13780 5731
rect 13722 5706 13758 5723
rect 13775 5706 13780 5723
rect 13722 5689 13780 5706
rect 13722 5672 13758 5689
rect 13775 5672 13780 5689
rect 13722 5655 13780 5672
rect 13722 5638 13758 5655
rect 13775 5638 13780 5655
rect 13722 5630 13780 5638
rect 13797 5723 13824 5731
rect 13797 5706 13802 5723
rect 13819 5706 13824 5723
rect 13797 5689 13824 5706
rect 13797 5672 13802 5689
rect 13819 5672 13824 5689
rect 13797 5655 13824 5672
rect 13797 5638 13802 5655
rect 13819 5638 13824 5655
rect 13186 5596 13190 5615
rect 13209 5596 13213 5615
rect 13797 5615 13824 5638
rect 13841 5723 13899 5731
rect 13841 5706 13846 5723
rect 13863 5706 13899 5723
rect 13841 5689 13899 5706
rect 13841 5672 13846 5689
rect 13863 5672 13899 5689
rect 13841 5655 13899 5672
rect 13841 5638 13846 5655
rect 13863 5638 13899 5655
rect 13841 5630 13899 5638
rect 13921 5723 13948 5731
rect 13921 5706 13926 5723
rect 13943 5706 13948 5723
rect 13921 5689 13948 5706
rect 13921 5672 13926 5689
rect 13943 5672 13948 5689
rect 13921 5655 13948 5672
rect 13921 5638 13926 5655
rect 13943 5638 13948 5655
rect 13921 5630 13948 5638
rect 14251 5723 14278 5731
rect 14251 5706 14256 5723
rect 14273 5706 14278 5723
rect 14251 5689 14278 5706
rect 14251 5672 14256 5689
rect 14273 5672 14278 5689
rect 14251 5655 14278 5672
rect 14251 5638 14256 5655
rect 14273 5638 14278 5655
rect 14251 5630 14278 5638
rect 14300 5723 14358 5731
rect 14300 5706 14336 5723
rect 14353 5706 14358 5723
rect 14300 5689 14358 5706
rect 14300 5672 14336 5689
rect 14353 5672 14358 5689
rect 14300 5655 14358 5672
rect 14300 5638 14336 5655
rect 14353 5638 14358 5655
rect 14300 5630 14358 5638
rect 14375 5723 14402 5731
rect 14375 5706 14380 5723
rect 14397 5706 14402 5723
rect 14375 5689 14402 5706
rect 14375 5672 14380 5689
rect 14397 5672 14402 5689
rect 14375 5655 14402 5672
rect 14375 5638 14380 5655
rect 14397 5638 14402 5655
rect 13797 5596 13801 5615
rect 13820 5596 13824 5615
rect 14375 5615 14402 5638
rect 14419 5723 14477 5731
rect 14419 5706 14424 5723
rect 14441 5706 14477 5723
rect 14419 5689 14477 5706
rect 14419 5672 14424 5689
rect 14441 5672 14477 5689
rect 14419 5655 14477 5672
rect 14419 5638 14424 5655
rect 14441 5638 14477 5655
rect 14419 5630 14477 5638
rect 14499 5723 14526 5731
rect 14499 5706 14504 5723
rect 14521 5706 14526 5723
rect 14499 5689 14526 5706
rect 14499 5672 14504 5689
rect 14521 5672 14526 5689
rect 14499 5655 14526 5672
rect 14499 5638 14504 5655
rect 14521 5638 14526 5655
rect 14499 5630 14526 5638
rect 14862 5723 14889 5731
rect 14862 5706 14867 5723
rect 14884 5706 14889 5723
rect 14862 5689 14889 5706
rect 14862 5672 14867 5689
rect 14884 5672 14889 5689
rect 14862 5655 14889 5672
rect 14862 5638 14867 5655
rect 14884 5638 14889 5655
rect 14862 5630 14889 5638
rect 14911 5723 14969 5731
rect 14911 5706 14947 5723
rect 14964 5706 14969 5723
rect 14911 5689 14969 5706
rect 14911 5672 14947 5689
rect 14964 5672 14969 5689
rect 14911 5655 14969 5672
rect 14911 5638 14947 5655
rect 14964 5638 14969 5655
rect 14911 5630 14969 5638
rect 14986 5723 15013 5731
rect 14986 5706 14991 5723
rect 15008 5706 15013 5723
rect 14986 5689 15013 5706
rect 14986 5672 14991 5689
rect 15008 5672 15013 5689
rect 14986 5655 15013 5672
rect 14986 5638 14991 5655
rect 15008 5638 15013 5655
rect 14375 5596 14379 5615
rect 14398 5596 14402 5615
rect 14986 5615 15013 5638
rect 15030 5723 15088 5731
rect 15030 5706 15035 5723
rect 15052 5706 15088 5723
rect 15030 5689 15088 5706
rect 15030 5672 15035 5689
rect 15052 5672 15088 5689
rect 15030 5655 15088 5672
rect 15030 5638 15035 5655
rect 15052 5638 15088 5655
rect 15030 5630 15088 5638
rect 15110 5723 15137 5731
rect 15110 5706 15115 5723
rect 15132 5706 15137 5723
rect 15110 5689 15137 5706
rect 15110 5672 15115 5689
rect 15132 5672 15137 5689
rect 15110 5655 15137 5672
rect 15110 5638 15115 5655
rect 15132 5638 15137 5655
rect 15110 5630 15137 5638
rect 15473 5723 15500 5731
rect 15473 5706 15478 5723
rect 15495 5706 15500 5723
rect 15473 5689 15500 5706
rect 15473 5672 15478 5689
rect 15495 5672 15500 5689
rect 15473 5655 15500 5672
rect 15473 5638 15478 5655
rect 15495 5638 15500 5655
rect 15473 5630 15500 5638
rect 15522 5723 15580 5731
rect 15522 5706 15558 5723
rect 15575 5706 15580 5723
rect 15522 5689 15580 5706
rect 15522 5672 15558 5689
rect 15575 5672 15580 5689
rect 15522 5655 15580 5672
rect 15522 5638 15558 5655
rect 15575 5638 15580 5655
rect 15522 5630 15580 5638
rect 15597 5723 15624 5731
rect 15597 5706 15602 5723
rect 15619 5706 15624 5723
rect 15597 5689 15624 5706
rect 15597 5672 15602 5689
rect 15619 5672 15624 5689
rect 15597 5655 15624 5672
rect 15597 5638 15602 5655
rect 15619 5638 15624 5655
rect 14986 5596 14990 5615
rect 15009 5596 15013 5615
rect 15597 5615 15624 5638
rect 15641 5723 15699 5731
rect 15641 5706 15646 5723
rect 15663 5706 15699 5723
rect 15641 5689 15699 5706
rect 15641 5672 15646 5689
rect 15663 5672 15699 5689
rect 15641 5655 15699 5672
rect 15641 5638 15646 5655
rect 15663 5638 15699 5655
rect 15641 5630 15699 5638
rect 15721 5723 15748 5731
rect 15721 5706 15726 5723
rect 15743 5706 15748 5723
rect 15721 5689 15748 5706
rect 15721 5672 15726 5689
rect 15743 5672 15748 5689
rect 15721 5655 15748 5672
rect 15721 5638 15726 5655
rect 15743 5638 15748 5655
rect 15721 5630 15748 5638
rect 15597 5596 15601 5615
rect 15620 5596 15624 5615
rect 12575 5472 12579 5491
rect 12598 5472 12602 5491
rect 12500 5449 12558 5457
rect 12500 5432 12536 5449
rect 12553 5432 12558 5449
rect 12500 5415 12558 5432
rect 12500 5398 12536 5415
rect 12553 5398 12558 5415
rect 12500 5381 12558 5398
rect 12500 5364 12536 5381
rect 12553 5364 12558 5381
rect 12500 5347 12558 5364
rect 12500 5330 12536 5347
rect 12553 5330 12558 5347
rect 12500 5313 12558 5330
rect 12500 5296 12536 5313
rect 12553 5296 12558 5313
rect 12500 5279 12558 5296
rect 12500 5262 12536 5279
rect 12553 5262 12558 5279
rect 12500 5254 12558 5262
rect 12575 5449 12602 5472
rect 13186 5472 13190 5491
rect 13209 5472 13213 5491
rect 12575 5432 12580 5449
rect 12597 5432 12602 5449
rect 12575 5415 12602 5432
rect 12575 5398 12580 5415
rect 12597 5398 12602 5415
rect 12575 5381 12602 5398
rect 12575 5364 12580 5381
rect 12597 5364 12602 5381
rect 12575 5347 12602 5364
rect 12575 5330 12580 5347
rect 12597 5330 12602 5347
rect 12575 5313 12602 5330
rect 12575 5296 12580 5313
rect 12597 5296 12602 5313
rect 12575 5279 12602 5296
rect 12575 5262 12580 5279
rect 12597 5262 12602 5279
rect 12575 5254 12602 5262
rect 12619 5449 12677 5457
rect 12619 5432 12624 5449
rect 12641 5432 12677 5449
rect 12619 5415 12677 5432
rect 12619 5398 12624 5415
rect 12641 5398 12677 5415
rect 12619 5381 12677 5398
rect 12619 5364 12624 5381
rect 12641 5364 12677 5381
rect 12619 5347 12677 5364
rect 12619 5330 12624 5347
rect 12641 5330 12677 5347
rect 12619 5313 12677 5330
rect 12619 5296 12624 5313
rect 12641 5296 12677 5313
rect 12619 5279 12677 5296
rect 12619 5262 12624 5279
rect 12641 5262 12677 5279
rect 12619 5254 12677 5262
rect 12450 5177 12483 5185
rect 12450 5160 12458 5177
rect 12475 5160 12483 5177
rect 12450 5152 12483 5160
rect 12500 5167 12527 5254
rect 12549 5229 12582 5237
rect 12549 5212 12557 5229
rect 12574 5221 12582 5229
rect 12650 5221 12677 5254
rect 12574 5212 12677 5221
rect 12549 5204 12677 5212
rect 12595 5175 12628 5183
rect 12595 5167 12603 5175
rect 12500 5158 12603 5167
rect 12620 5158 12628 5175
rect 12500 5150 12628 5158
rect 12450 5123 12483 5131
rect 12450 5106 12458 5123
rect 12475 5106 12483 5123
rect 12450 5098 12483 5106
rect 12500 5081 12527 5150
rect 12650 5081 12677 5204
rect 13111 5449 13169 5457
rect 13111 5432 13147 5449
rect 13164 5432 13169 5449
rect 13111 5415 13169 5432
rect 13111 5398 13147 5415
rect 13164 5398 13169 5415
rect 13111 5381 13169 5398
rect 13111 5364 13147 5381
rect 13164 5364 13169 5381
rect 13111 5347 13169 5364
rect 13111 5330 13147 5347
rect 13164 5330 13169 5347
rect 13111 5313 13169 5330
rect 13111 5296 13147 5313
rect 13164 5296 13169 5313
rect 13111 5279 13169 5296
rect 13111 5262 13147 5279
rect 13164 5262 13169 5279
rect 13111 5254 13169 5262
rect 13186 5449 13213 5472
rect 13797 5472 13801 5491
rect 13820 5472 13824 5491
rect 13186 5432 13191 5449
rect 13208 5432 13213 5449
rect 13186 5415 13213 5432
rect 13186 5398 13191 5415
rect 13208 5398 13213 5415
rect 13186 5381 13213 5398
rect 13186 5364 13191 5381
rect 13208 5364 13213 5381
rect 13186 5347 13213 5364
rect 13186 5330 13191 5347
rect 13208 5330 13213 5347
rect 13186 5313 13213 5330
rect 13186 5296 13191 5313
rect 13208 5296 13213 5313
rect 13186 5279 13213 5296
rect 13186 5262 13191 5279
rect 13208 5262 13213 5279
rect 13186 5254 13213 5262
rect 13230 5449 13288 5457
rect 13230 5432 13235 5449
rect 13252 5432 13288 5449
rect 13230 5415 13288 5432
rect 13230 5398 13235 5415
rect 13252 5398 13288 5415
rect 13230 5381 13288 5398
rect 13230 5364 13235 5381
rect 13252 5364 13288 5381
rect 13230 5347 13288 5364
rect 13230 5330 13235 5347
rect 13252 5330 13288 5347
rect 13230 5313 13288 5330
rect 13230 5296 13235 5313
rect 13252 5296 13288 5313
rect 13230 5279 13288 5296
rect 13230 5262 13235 5279
rect 13252 5262 13288 5279
rect 13230 5254 13288 5262
rect 13061 5177 13094 5185
rect 13061 5160 13069 5177
rect 13086 5160 13094 5177
rect 13061 5152 13094 5160
rect 13111 5167 13138 5254
rect 13160 5229 13193 5237
rect 13160 5212 13168 5229
rect 13185 5221 13193 5229
rect 13261 5221 13288 5254
rect 13185 5212 13288 5221
rect 13160 5204 13288 5212
rect 13206 5175 13239 5183
rect 13206 5167 13214 5175
rect 13111 5158 13214 5167
rect 13231 5158 13239 5175
rect 13111 5150 13239 5158
rect 12694 5139 12727 5147
rect 12694 5122 12702 5139
rect 12719 5122 12727 5139
rect 12694 5114 12727 5122
rect 13061 5123 13094 5131
rect 13061 5106 13069 5123
rect 13086 5106 13094 5123
rect 13061 5098 13094 5106
rect 13111 5081 13138 5150
rect 13261 5081 13288 5204
rect 13722 5449 13780 5457
rect 13722 5432 13758 5449
rect 13775 5432 13780 5449
rect 13722 5415 13780 5432
rect 13722 5398 13758 5415
rect 13775 5398 13780 5415
rect 13722 5381 13780 5398
rect 13722 5364 13758 5381
rect 13775 5364 13780 5381
rect 13722 5347 13780 5364
rect 13722 5330 13758 5347
rect 13775 5330 13780 5347
rect 13722 5313 13780 5330
rect 13722 5296 13758 5313
rect 13775 5296 13780 5313
rect 13722 5279 13780 5296
rect 13722 5262 13758 5279
rect 13775 5262 13780 5279
rect 13722 5254 13780 5262
rect 13797 5449 13824 5472
rect 14375 5472 14379 5491
rect 14398 5472 14402 5491
rect 13797 5432 13802 5449
rect 13819 5432 13824 5449
rect 13797 5415 13824 5432
rect 13797 5398 13802 5415
rect 13819 5398 13824 5415
rect 13797 5381 13824 5398
rect 13797 5364 13802 5381
rect 13819 5364 13824 5381
rect 13797 5347 13824 5364
rect 13797 5330 13802 5347
rect 13819 5330 13824 5347
rect 13797 5313 13824 5330
rect 13797 5296 13802 5313
rect 13819 5296 13824 5313
rect 13797 5279 13824 5296
rect 13797 5262 13802 5279
rect 13819 5262 13824 5279
rect 13797 5254 13824 5262
rect 13841 5449 13899 5457
rect 13841 5432 13846 5449
rect 13863 5432 13899 5449
rect 13841 5415 13899 5432
rect 13841 5398 13846 5415
rect 13863 5398 13899 5415
rect 13841 5381 13899 5398
rect 13841 5364 13846 5381
rect 13863 5364 13899 5381
rect 13841 5347 13899 5364
rect 13841 5330 13846 5347
rect 13863 5330 13899 5347
rect 13841 5313 13899 5330
rect 13841 5296 13846 5313
rect 13863 5296 13899 5313
rect 13841 5279 13899 5296
rect 13841 5262 13846 5279
rect 13863 5262 13899 5279
rect 13841 5254 13899 5262
rect 13672 5177 13705 5185
rect 13672 5160 13680 5177
rect 13697 5160 13705 5177
rect 13672 5152 13705 5160
rect 13722 5167 13749 5254
rect 13771 5229 13804 5237
rect 13771 5212 13779 5229
rect 13796 5221 13804 5229
rect 13872 5221 13899 5254
rect 13796 5212 13899 5221
rect 13771 5204 13899 5212
rect 13817 5175 13850 5183
rect 13817 5167 13825 5175
rect 13722 5158 13825 5167
rect 13842 5158 13850 5175
rect 13722 5150 13850 5158
rect 13305 5139 13338 5147
rect 13305 5122 13313 5139
rect 13330 5122 13338 5139
rect 13305 5114 13338 5122
rect 13672 5123 13705 5131
rect 13672 5106 13680 5123
rect 13697 5106 13705 5123
rect 13672 5098 13705 5106
rect 13722 5081 13749 5150
rect 13872 5081 13899 5204
rect 14300 5449 14358 5457
rect 14300 5432 14336 5449
rect 14353 5432 14358 5449
rect 14300 5415 14358 5432
rect 14300 5398 14336 5415
rect 14353 5398 14358 5415
rect 14300 5381 14358 5398
rect 14300 5364 14336 5381
rect 14353 5364 14358 5381
rect 14300 5347 14358 5364
rect 14300 5330 14336 5347
rect 14353 5330 14358 5347
rect 14300 5313 14358 5330
rect 14300 5296 14336 5313
rect 14353 5296 14358 5313
rect 14300 5279 14358 5296
rect 14300 5262 14336 5279
rect 14353 5262 14358 5279
rect 14300 5254 14358 5262
rect 14375 5449 14402 5472
rect 14986 5472 14990 5491
rect 15009 5472 15013 5491
rect 14375 5432 14380 5449
rect 14397 5432 14402 5449
rect 14375 5415 14402 5432
rect 14375 5398 14380 5415
rect 14397 5398 14402 5415
rect 14375 5381 14402 5398
rect 14375 5364 14380 5381
rect 14397 5364 14402 5381
rect 14375 5347 14402 5364
rect 14375 5330 14380 5347
rect 14397 5330 14402 5347
rect 14375 5313 14402 5330
rect 14375 5296 14380 5313
rect 14397 5296 14402 5313
rect 14375 5279 14402 5296
rect 14375 5262 14380 5279
rect 14397 5262 14402 5279
rect 14375 5254 14402 5262
rect 14419 5449 14477 5457
rect 14419 5432 14424 5449
rect 14441 5432 14477 5449
rect 14419 5415 14477 5432
rect 14419 5398 14424 5415
rect 14441 5398 14477 5415
rect 14419 5381 14477 5398
rect 14419 5364 14424 5381
rect 14441 5364 14477 5381
rect 14419 5347 14477 5364
rect 14419 5330 14424 5347
rect 14441 5330 14477 5347
rect 14419 5313 14477 5330
rect 14419 5296 14424 5313
rect 14441 5296 14477 5313
rect 14419 5279 14477 5296
rect 14419 5262 14424 5279
rect 14441 5262 14477 5279
rect 14419 5254 14477 5262
rect 14250 5177 14283 5185
rect 14250 5160 14258 5177
rect 14275 5160 14283 5177
rect 14250 5152 14283 5160
rect 14300 5167 14327 5254
rect 14349 5229 14382 5237
rect 14349 5212 14357 5229
rect 14374 5221 14382 5229
rect 14450 5221 14477 5254
rect 14374 5212 14477 5221
rect 14349 5204 14477 5212
rect 14395 5175 14428 5183
rect 14395 5167 14403 5175
rect 14300 5158 14403 5167
rect 14420 5158 14428 5175
rect 14300 5150 14428 5158
rect 13916 5139 13949 5147
rect 13916 5122 13924 5139
rect 13941 5122 13949 5139
rect 13916 5114 13949 5122
rect 14250 5123 14283 5131
rect 14250 5106 14258 5123
rect 14275 5106 14283 5123
rect 14250 5098 14283 5106
rect 14300 5081 14327 5150
rect 14450 5081 14477 5204
rect 14911 5449 14969 5457
rect 14911 5432 14947 5449
rect 14964 5432 14969 5449
rect 14911 5415 14969 5432
rect 14911 5398 14947 5415
rect 14964 5398 14969 5415
rect 14911 5381 14969 5398
rect 14911 5364 14947 5381
rect 14964 5364 14969 5381
rect 14911 5347 14969 5364
rect 14911 5330 14947 5347
rect 14964 5330 14969 5347
rect 14911 5313 14969 5330
rect 14911 5296 14947 5313
rect 14964 5296 14969 5313
rect 14911 5279 14969 5296
rect 14911 5262 14947 5279
rect 14964 5262 14969 5279
rect 14911 5254 14969 5262
rect 14986 5449 15013 5472
rect 15597 5472 15601 5491
rect 15620 5472 15624 5491
rect 14986 5432 14991 5449
rect 15008 5432 15013 5449
rect 14986 5415 15013 5432
rect 14986 5398 14991 5415
rect 15008 5398 15013 5415
rect 14986 5381 15013 5398
rect 14986 5364 14991 5381
rect 15008 5364 15013 5381
rect 14986 5347 15013 5364
rect 14986 5330 14991 5347
rect 15008 5330 15013 5347
rect 14986 5313 15013 5330
rect 14986 5296 14991 5313
rect 15008 5296 15013 5313
rect 14986 5279 15013 5296
rect 14986 5262 14991 5279
rect 15008 5262 15013 5279
rect 14986 5254 15013 5262
rect 15030 5449 15088 5457
rect 15030 5432 15035 5449
rect 15052 5432 15088 5449
rect 15030 5415 15088 5432
rect 15030 5398 15035 5415
rect 15052 5398 15088 5415
rect 15030 5381 15088 5398
rect 15030 5364 15035 5381
rect 15052 5364 15088 5381
rect 15030 5347 15088 5364
rect 15030 5330 15035 5347
rect 15052 5330 15088 5347
rect 15030 5313 15088 5330
rect 15030 5296 15035 5313
rect 15052 5296 15088 5313
rect 15030 5279 15088 5296
rect 15030 5262 15035 5279
rect 15052 5262 15088 5279
rect 15030 5254 15088 5262
rect 14861 5177 14894 5185
rect 14861 5160 14869 5177
rect 14886 5160 14894 5177
rect 14861 5152 14894 5160
rect 14911 5167 14938 5254
rect 14960 5229 14993 5237
rect 14960 5212 14968 5229
rect 14985 5221 14993 5229
rect 15061 5221 15088 5254
rect 14985 5212 15088 5221
rect 14960 5204 15088 5212
rect 15006 5175 15039 5183
rect 15006 5167 15014 5175
rect 14911 5158 15014 5167
rect 15031 5158 15039 5175
rect 14911 5150 15039 5158
rect 14494 5139 14527 5147
rect 14494 5122 14502 5139
rect 14519 5122 14527 5139
rect 14494 5114 14527 5122
rect 14861 5123 14894 5131
rect 14861 5106 14869 5123
rect 14886 5106 14894 5123
rect 14861 5098 14894 5106
rect 14911 5081 14938 5150
rect 15061 5081 15088 5204
rect 15522 5449 15580 5457
rect 15522 5432 15558 5449
rect 15575 5432 15580 5449
rect 15522 5415 15580 5432
rect 15522 5398 15558 5415
rect 15575 5398 15580 5415
rect 15522 5381 15580 5398
rect 15522 5364 15558 5381
rect 15575 5364 15580 5381
rect 15522 5347 15580 5364
rect 15522 5330 15558 5347
rect 15575 5330 15580 5347
rect 15522 5313 15580 5330
rect 15522 5296 15558 5313
rect 15575 5296 15580 5313
rect 15522 5279 15580 5296
rect 15522 5262 15558 5279
rect 15575 5262 15580 5279
rect 15522 5254 15580 5262
rect 15597 5449 15624 5472
rect 15597 5432 15602 5449
rect 15619 5432 15624 5449
rect 15597 5415 15624 5432
rect 15597 5398 15602 5415
rect 15619 5398 15624 5415
rect 15597 5381 15624 5398
rect 15597 5364 15602 5381
rect 15619 5364 15624 5381
rect 15597 5347 15624 5364
rect 15597 5330 15602 5347
rect 15619 5330 15624 5347
rect 15597 5313 15624 5330
rect 15597 5296 15602 5313
rect 15619 5296 15624 5313
rect 15597 5279 15624 5296
rect 15597 5262 15602 5279
rect 15619 5262 15624 5279
rect 15597 5254 15624 5262
rect 15641 5449 15699 5457
rect 15641 5432 15646 5449
rect 15663 5432 15699 5449
rect 15641 5415 15699 5432
rect 15641 5398 15646 5415
rect 15663 5398 15699 5415
rect 15641 5381 15699 5398
rect 15641 5364 15646 5381
rect 15663 5364 15699 5381
rect 15641 5347 15699 5364
rect 15641 5330 15646 5347
rect 15663 5330 15699 5347
rect 15641 5313 15699 5330
rect 15641 5296 15646 5313
rect 15663 5296 15699 5313
rect 15641 5279 15699 5296
rect 15641 5262 15646 5279
rect 15663 5262 15699 5279
rect 15641 5254 15699 5262
rect 15472 5177 15505 5185
rect 15472 5160 15480 5177
rect 15497 5160 15505 5177
rect 15472 5152 15505 5160
rect 15522 5167 15549 5254
rect 15571 5229 15604 5237
rect 15571 5212 15579 5229
rect 15596 5221 15604 5229
rect 15672 5221 15699 5254
rect 15596 5212 15699 5221
rect 15571 5204 15699 5212
rect 15617 5175 15650 5183
rect 15617 5167 15625 5175
rect 15522 5158 15625 5167
rect 15642 5158 15650 5175
rect 15522 5150 15650 5158
rect 15105 5139 15138 5147
rect 15105 5122 15113 5139
rect 15130 5122 15138 5139
rect 15105 5114 15138 5122
rect 15472 5123 15505 5131
rect 15472 5106 15480 5123
rect 15497 5106 15505 5123
rect 15472 5098 15505 5106
rect 15522 5081 15549 5150
rect 15672 5081 15699 5204
rect 15716 5139 15749 5147
rect 15716 5122 15724 5139
rect 15741 5122 15749 5139
rect 15716 5114 15749 5122
rect 12451 5073 12478 5081
rect 12451 5056 12456 5073
rect 12473 5056 12478 5073
rect 12451 5039 12478 5056
rect 12451 5022 12456 5039
rect 12473 5022 12478 5039
rect 12451 5005 12478 5022
rect 12451 4988 12456 5005
rect 12473 4988 12478 5005
rect 12451 4980 12478 4988
rect 12500 5073 12558 5081
rect 12500 5056 12536 5073
rect 12553 5056 12558 5073
rect 12500 5039 12558 5056
rect 12500 5022 12536 5039
rect 12553 5022 12558 5039
rect 12500 5005 12558 5022
rect 12500 4988 12536 5005
rect 12553 4988 12558 5005
rect 12500 4980 12558 4988
rect 12575 5073 12602 5081
rect 12575 5056 12580 5073
rect 12597 5056 12602 5073
rect 12575 5039 12602 5056
rect 12575 5022 12580 5039
rect 12597 5022 12602 5039
rect 12575 5005 12602 5022
rect 12575 4988 12580 5005
rect 12597 4988 12602 5005
rect 12575 4965 12602 4988
rect 12619 5073 12677 5081
rect 12619 5056 12624 5073
rect 12641 5056 12677 5073
rect 12619 5039 12677 5056
rect 12619 5022 12624 5039
rect 12641 5022 12677 5039
rect 12619 5005 12677 5022
rect 12619 4988 12624 5005
rect 12641 4988 12677 5005
rect 12619 4980 12677 4988
rect 12699 5073 12726 5081
rect 12699 5056 12704 5073
rect 12721 5056 12726 5073
rect 12699 5039 12726 5056
rect 12699 5022 12704 5039
rect 12721 5022 12726 5039
rect 12699 5005 12726 5022
rect 12699 4988 12704 5005
rect 12721 4988 12726 5005
rect 12699 4980 12726 4988
rect 13062 5073 13089 5081
rect 13062 5056 13067 5073
rect 13084 5056 13089 5073
rect 13062 5039 13089 5056
rect 13062 5022 13067 5039
rect 13084 5022 13089 5039
rect 13062 5005 13089 5022
rect 13062 4988 13067 5005
rect 13084 4988 13089 5005
rect 13062 4980 13089 4988
rect 13111 5073 13169 5081
rect 13111 5056 13147 5073
rect 13164 5056 13169 5073
rect 13111 5039 13169 5056
rect 13111 5022 13147 5039
rect 13164 5022 13169 5039
rect 13111 5005 13169 5022
rect 13111 4988 13147 5005
rect 13164 4988 13169 5005
rect 13111 4980 13169 4988
rect 13186 5073 13213 5081
rect 13186 5056 13191 5073
rect 13208 5056 13213 5073
rect 13186 5039 13213 5056
rect 13186 5022 13191 5039
rect 13208 5022 13213 5039
rect 13186 5005 13213 5022
rect 13186 4988 13191 5005
rect 13208 4988 13213 5005
rect 12575 4946 12579 4965
rect 12598 4946 12602 4965
rect 13186 4965 13213 4988
rect 13230 5073 13288 5081
rect 13230 5056 13235 5073
rect 13252 5056 13288 5073
rect 13230 5039 13288 5056
rect 13230 5022 13235 5039
rect 13252 5022 13288 5039
rect 13230 5005 13288 5022
rect 13230 4988 13235 5005
rect 13252 4988 13288 5005
rect 13230 4980 13288 4988
rect 13310 5073 13337 5081
rect 13310 5056 13315 5073
rect 13332 5056 13337 5073
rect 13310 5039 13337 5056
rect 13310 5022 13315 5039
rect 13332 5022 13337 5039
rect 13310 5005 13337 5022
rect 13310 4988 13315 5005
rect 13332 4988 13337 5005
rect 13310 4980 13337 4988
rect 13673 5073 13700 5081
rect 13673 5056 13678 5073
rect 13695 5056 13700 5073
rect 13673 5039 13700 5056
rect 13673 5022 13678 5039
rect 13695 5022 13700 5039
rect 13673 5005 13700 5022
rect 13673 4988 13678 5005
rect 13695 4988 13700 5005
rect 13673 4980 13700 4988
rect 13722 5073 13780 5081
rect 13722 5056 13758 5073
rect 13775 5056 13780 5073
rect 13722 5039 13780 5056
rect 13722 5022 13758 5039
rect 13775 5022 13780 5039
rect 13722 5005 13780 5022
rect 13722 4988 13758 5005
rect 13775 4988 13780 5005
rect 13722 4980 13780 4988
rect 13797 5073 13824 5081
rect 13797 5056 13802 5073
rect 13819 5056 13824 5073
rect 13797 5039 13824 5056
rect 13797 5022 13802 5039
rect 13819 5022 13824 5039
rect 13797 5005 13824 5022
rect 13797 4988 13802 5005
rect 13819 4988 13824 5005
rect 13186 4946 13190 4965
rect 13209 4946 13213 4965
rect 13797 4965 13824 4988
rect 13841 5073 13899 5081
rect 13841 5056 13846 5073
rect 13863 5056 13899 5073
rect 13841 5039 13899 5056
rect 13841 5022 13846 5039
rect 13863 5022 13899 5039
rect 13841 5005 13899 5022
rect 13841 4988 13846 5005
rect 13863 4988 13899 5005
rect 13841 4980 13899 4988
rect 13921 5073 13948 5081
rect 13921 5056 13926 5073
rect 13943 5056 13948 5073
rect 13921 5039 13948 5056
rect 13921 5022 13926 5039
rect 13943 5022 13948 5039
rect 13921 5005 13948 5022
rect 13921 4988 13926 5005
rect 13943 4988 13948 5005
rect 13921 4980 13948 4988
rect 14251 5073 14278 5081
rect 14251 5056 14256 5073
rect 14273 5056 14278 5073
rect 14251 5039 14278 5056
rect 14251 5022 14256 5039
rect 14273 5022 14278 5039
rect 14251 5005 14278 5022
rect 14251 4988 14256 5005
rect 14273 4988 14278 5005
rect 14251 4980 14278 4988
rect 14300 5073 14358 5081
rect 14300 5056 14336 5073
rect 14353 5056 14358 5073
rect 14300 5039 14358 5056
rect 14300 5022 14336 5039
rect 14353 5022 14358 5039
rect 14300 5005 14358 5022
rect 14300 4988 14336 5005
rect 14353 4988 14358 5005
rect 14300 4980 14358 4988
rect 14375 5073 14402 5081
rect 14375 5056 14380 5073
rect 14397 5056 14402 5073
rect 14375 5039 14402 5056
rect 14375 5022 14380 5039
rect 14397 5022 14402 5039
rect 14375 5005 14402 5022
rect 14375 4988 14380 5005
rect 14397 4988 14402 5005
rect 13797 4946 13801 4965
rect 13820 4946 13824 4965
rect 14375 4965 14402 4988
rect 14419 5073 14477 5081
rect 14419 5056 14424 5073
rect 14441 5056 14477 5073
rect 14419 5039 14477 5056
rect 14419 5022 14424 5039
rect 14441 5022 14477 5039
rect 14419 5005 14477 5022
rect 14419 4988 14424 5005
rect 14441 4988 14477 5005
rect 14419 4980 14477 4988
rect 14499 5073 14526 5081
rect 14499 5056 14504 5073
rect 14521 5056 14526 5073
rect 14499 5039 14526 5056
rect 14499 5022 14504 5039
rect 14521 5022 14526 5039
rect 14499 5005 14526 5022
rect 14499 4988 14504 5005
rect 14521 4988 14526 5005
rect 14499 4980 14526 4988
rect 14862 5073 14889 5081
rect 14862 5056 14867 5073
rect 14884 5056 14889 5073
rect 14862 5039 14889 5056
rect 14862 5022 14867 5039
rect 14884 5022 14889 5039
rect 14862 5005 14889 5022
rect 14862 4988 14867 5005
rect 14884 4988 14889 5005
rect 14862 4980 14889 4988
rect 14911 5073 14969 5081
rect 14911 5056 14947 5073
rect 14964 5056 14969 5073
rect 14911 5039 14969 5056
rect 14911 5022 14947 5039
rect 14964 5022 14969 5039
rect 14911 5005 14969 5022
rect 14911 4988 14947 5005
rect 14964 4988 14969 5005
rect 14911 4980 14969 4988
rect 14986 5073 15013 5081
rect 14986 5056 14991 5073
rect 15008 5056 15013 5073
rect 14986 5039 15013 5056
rect 14986 5022 14991 5039
rect 15008 5022 15013 5039
rect 14986 5005 15013 5022
rect 14986 4988 14991 5005
rect 15008 4988 15013 5005
rect 14375 4946 14379 4965
rect 14398 4946 14402 4965
rect 14986 4965 15013 4988
rect 15030 5073 15088 5081
rect 15030 5056 15035 5073
rect 15052 5056 15088 5073
rect 15030 5039 15088 5056
rect 15030 5022 15035 5039
rect 15052 5022 15088 5039
rect 15030 5005 15088 5022
rect 15030 4988 15035 5005
rect 15052 4988 15088 5005
rect 15030 4980 15088 4988
rect 15110 5073 15137 5081
rect 15110 5056 15115 5073
rect 15132 5056 15137 5073
rect 15110 5039 15137 5056
rect 15110 5022 15115 5039
rect 15132 5022 15137 5039
rect 15110 5005 15137 5022
rect 15110 4988 15115 5005
rect 15132 4988 15137 5005
rect 15110 4980 15137 4988
rect 15473 5073 15500 5081
rect 15473 5056 15478 5073
rect 15495 5056 15500 5073
rect 15473 5039 15500 5056
rect 15473 5022 15478 5039
rect 15495 5022 15500 5039
rect 15473 5005 15500 5022
rect 15473 4988 15478 5005
rect 15495 4988 15500 5005
rect 15473 4980 15500 4988
rect 15522 5073 15580 5081
rect 15522 5056 15558 5073
rect 15575 5056 15580 5073
rect 15522 5039 15580 5056
rect 15522 5022 15558 5039
rect 15575 5022 15580 5039
rect 15522 5005 15580 5022
rect 15522 4988 15558 5005
rect 15575 4988 15580 5005
rect 15522 4980 15580 4988
rect 15597 5073 15624 5081
rect 15597 5056 15602 5073
rect 15619 5056 15624 5073
rect 15597 5039 15624 5056
rect 15597 5022 15602 5039
rect 15619 5022 15624 5039
rect 15597 5005 15624 5022
rect 15597 4988 15602 5005
rect 15619 4988 15624 5005
rect 14986 4946 14990 4965
rect 15009 4946 15013 4965
rect 15597 4965 15624 4988
rect 15641 5073 15699 5081
rect 15641 5056 15646 5073
rect 15663 5056 15699 5073
rect 15641 5039 15699 5056
rect 15641 5022 15646 5039
rect 15663 5022 15699 5039
rect 15641 5005 15699 5022
rect 15641 4988 15646 5005
rect 15663 4988 15699 5005
rect 15641 4980 15699 4988
rect 15721 5073 15748 5081
rect 15721 5056 15726 5073
rect 15743 5056 15748 5073
rect 15721 5039 15748 5056
rect 15721 5022 15726 5039
rect 15743 5022 15748 5039
rect 15721 5005 15748 5022
rect 15721 4988 15726 5005
rect 15743 4988 15748 5005
rect 15721 4980 15748 4988
rect 15597 4946 15601 4965
rect 15620 4946 15624 4965
rect 12575 4832 12579 4851
rect 12598 4832 12602 4851
rect 12500 4809 12558 4817
rect 12500 4792 12536 4809
rect 12553 4792 12558 4809
rect 12500 4775 12558 4792
rect 12500 4758 12536 4775
rect 12553 4758 12558 4775
rect 12500 4741 12558 4758
rect 12500 4724 12536 4741
rect 12553 4724 12558 4741
rect 12500 4707 12558 4724
rect 12500 4690 12536 4707
rect 12553 4690 12558 4707
rect 12500 4673 12558 4690
rect 12500 4656 12536 4673
rect 12553 4656 12558 4673
rect 12500 4639 12558 4656
rect 12500 4622 12536 4639
rect 12553 4622 12558 4639
rect 12500 4614 12558 4622
rect 12575 4809 12602 4832
rect 13186 4832 13190 4851
rect 13209 4832 13213 4851
rect 12575 4792 12580 4809
rect 12597 4792 12602 4809
rect 12575 4775 12602 4792
rect 12575 4758 12580 4775
rect 12597 4758 12602 4775
rect 12575 4741 12602 4758
rect 12575 4724 12580 4741
rect 12597 4724 12602 4741
rect 12575 4707 12602 4724
rect 12575 4690 12580 4707
rect 12597 4690 12602 4707
rect 12575 4673 12602 4690
rect 12575 4656 12580 4673
rect 12597 4656 12602 4673
rect 12575 4639 12602 4656
rect 12575 4622 12580 4639
rect 12597 4622 12602 4639
rect 12575 4614 12602 4622
rect 12619 4809 12677 4817
rect 12619 4792 12624 4809
rect 12641 4792 12677 4809
rect 12619 4775 12677 4792
rect 12619 4758 12624 4775
rect 12641 4758 12677 4775
rect 12619 4741 12677 4758
rect 12619 4724 12624 4741
rect 12641 4724 12677 4741
rect 12619 4707 12677 4724
rect 12619 4690 12624 4707
rect 12641 4690 12677 4707
rect 12619 4673 12677 4690
rect 12619 4656 12624 4673
rect 12641 4656 12677 4673
rect 12619 4639 12677 4656
rect 12619 4622 12624 4639
rect 12641 4622 12677 4639
rect 12619 4614 12677 4622
rect 12450 4537 12483 4545
rect 12450 4520 12458 4537
rect 12475 4520 12483 4537
rect 12450 4512 12483 4520
rect 12500 4527 12527 4614
rect 12549 4589 12582 4597
rect 12549 4572 12557 4589
rect 12574 4581 12582 4589
rect 12650 4581 12677 4614
rect 12574 4572 12677 4581
rect 12549 4564 12677 4572
rect 12595 4535 12628 4543
rect 12595 4527 12603 4535
rect 12500 4518 12603 4527
rect 12620 4518 12628 4535
rect 12500 4510 12628 4518
rect 12450 4483 12483 4491
rect 12450 4466 12458 4483
rect 12475 4466 12483 4483
rect 12450 4458 12483 4466
rect 12500 4441 12527 4510
rect 12650 4441 12677 4564
rect 13111 4809 13169 4817
rect 13111 4792 13147 4809
rect 13164 4792 13169 4809
rect 13111 4775 13169 4792
rect 13111 4758 13147 4775
rect 13164 4758 13169 4775
rect 13111 4741 13169 4758
rect 13111 4724 13147 4741
rect 13164 4724 13169 4741
rect 13111 4707 13169 4724
rect 13111 4690 13147 4707
rect 13164 4690 13169 4707
rect 13111 4673 13169 4690
rect 13111 4656 13147 4673
rect 13164 4656 13169 4673
rect 13111 4639 13169 4656
rect 13111 4622 13147 4639
rect 13164 4622 13169 4639
rect 13111 4614 13169 4622
rect 13186 4809 13213 4832
rect 13797 4832 13801 4851
rect 13820 4832 13824 4851
rect 13186 4792 13191 4809
rect 13208 4792 13213 4809
rect 13186 4775 13213 4792
rect 13186 4758 13191 4775
rect 13208 4758 13213 4775
rect 13186 4741 13213 4758
rect 13186 4724 13191 4741
rect 13208 4724 13213 4741
rect 13186 4707 13213 4724
rect 13186 4690 13191 4707
rect 13208 4690 13213 4707
rect 13186 4673 13213 4690
rect 13186 4656 13191 4673
rect 13208 4656 13213 4673
rect 13186 4639 13213 4656
rect 13186 4622 13191 4639
rect 13208 4622 13213 4639
rect 13186 4614 13213 4622
rect 13230 4809 13288 4817
rect 13230 4792 13235 4809
rect 13252 4792 13288 4809
rect 13230 4775 13288 4792
rect 13230 4758 13235 4775
rect 13252 4758 13288 4775
rect 13230 4741 13288 4758
rect 13230 4724 13235 4741
rect 13252 4724 13288 4741
rect 13230 4707 13288 4724
rect 13230 4690 13235 4707
rect 13252 4690 13288 4707
rect 13230 4673 13288 4690
rect 13230 4656 13235 4673
rect 13252 4656 13288 4673
rect 13230 4639 13288 4656
rect 13230 4622 13235 4639
rect 13252 4622 13288 4639
rect 13230 4614 13288 4622
rect 13061 4537 13094 4545
rect 13061 4520 13069 4537
rect 13086 4520 13094 4537
rect 13061 4512 13094 4520
rect 13111 4527 13138 4614
rect 13160 4589 13193 4597
rect 13160 4572 13168 4589
rect 13185 4581 13193 4589
rect 13261 4581 13288 4614
rect 13185 4572 13288 4581
rect 13160 4564 13288 4572
rect 13206 4535 13239 4543
rect 13206 4527 13214 4535
rect 13111 4518 13214 4527
rect 13231 4518 13239 4535
rect 13111 4510 13239 4518
rect 12694 4499 12727 4507
rect 12694 4482 12702 4499
rect 12719 4482 12727 4499
rect 12694 4474 12727 4482
rect 13061 4483 13094 4491
rect 13061 4466 13069 4483
rect 13086 4466 13094 4483
rect 13061 4458 13094 4466
rect 13111 4441 13138 4510
rect 13261 4441 13288 4564
rect 13722 4809 13780 4817
rect 13722 4792 13758 4809
rect 13775 4792 13780 4809
rect 13722 4775 13780 4792
rect 13722 4758 13758 4775
rect 13775 4758 13780 4775
rect 13722 4741 13780 4758
rect 13722 4724 13758 4741
rect 13775 4724 13780 4741
rect 13722 4707 13780 4724
rect 13722 4690 13758 4707
rect 13775 4690 13780 4707
rect 13722 4673 13780 4690
rect 13722 4656 13758 4673
rect 13775 4656 13780 4673
rect 13722 4639 13780 4656
rect 13722 4622 13758 4639
rect 13775 4622 13780 4639
rect 13722 4614 13780 4622
rect 13797 4809 13824 4832
rect 14375 4832 14379 4851
rect 14398 4832 14402 4851
rect 13797 4792 13802 4809
rect 13819 4792 13824 4809
rect 13797 4775 13824 4792
rect 13797 4758 13802 4775
rect 13819 4758 13824 4775
rect 13797 4741 13824 4758
rect 13797 4724 13802 4741
rect 13819 4724 13824 4741
rect 13797 4707 13824 4724
rect 13797 4690 13802 4707
rect 13819 4690 13824 4707
rect 13797 4673 13824 4690
rect 13797 4656 13802 4673
rect 13819 4656 13824 4673
rect 13797 4639 13824 4656
rect 13797 4622 13802 4639
rect 13819 4622 13824 4639
rect 13797 4614 13824 4622
rect 13841 4809 13899 4817
rect 13841 4792 13846 4809
rect 13863 4792 13899 4809
rect 13841 4775 13899 4792
rect 13841 4758 13846 4775
rect 13863 4758 13899 4775
rect 13841 4741 13899 4758
rect 13841 4724 13846 4741
rect 13863 4724 13899 4741
rect 13841 4707 13899 4724
rect 13841 4690 13846 4707
rect 13863 4690 13899 4707
rect 13841 4673 13899 4690
rect 13841 4656 13846 4673
rect 13863 4656 13899 4673
rect 13841 4639 13899 4656
rect 13841 4622 13846 4639
rect 13863 4622 13899 4639
rect 13841 4614 13899 4622
rect 13672 4537 13705 4545
rect 13672 4520 13680 4537
rect 13697 4520 13705 4537
rect 13672 4512 13705 4520
rect 13722 4527 13749 4614
rect 13771 4589 13804 4597
rect 13771 4572 13779 4589
rect 13796 4581 13804 4589
rect 13872 4581 13899 4614
rect 13796 4572 13899 4581
rect 13771 4564 13899 4572
rect 13817 4535 13850 4543
rect 13817 4527 13825 4535
rect 13722 4518 13825 4527
rect 13842 4518 13850 4535
rect 13722 4510 13850 4518
rect 13305 4499 13338 4507
rect 13305 4482 13313 4499
rect 13330 4482 13338 4499
rect 13305 4474 13338 4482
rect 13672 4483 13705 4491
rect 13672 4466 13680 4483
rect 13697 4466 13705 4483
rect 13672 4458 13705 4466
rect 13722 4441 13749 4510
rect 13872 4441 13899 4564
rect 14300 4809 14358 4817
rect 14300 4792 14336 4809
rect 14353 4792 14358 4809
rect 14300 4775 14358 4792
rect 14300 4758 14336 4775
rect 14353 4758 14358 4775
rect 14300 4741 14358 4758
rect 14300 4724 14336 4741
rect 14353 4724 14358 4741
rect 14300 4707 14358 4724
rect 14300 4690 14336 4707
rect 14353 4690 14358 4707
rect 14300 4673 14358 4690
rect 14300 4656 14336 4673
rect 14353 4656 14358 4673
rect 14300 4639 14358 4656
rect 14300 4622 14336 4639
rect 14353 4622 14358 4639
rect 14300 4614 14358 4622
rect 14375 4809 14402 4832
rect 14986 4832 14990 4851
rect 15009 4832 15013 4851
rect 14375 4792 14380 4809
rect 14397 4792 14402 4809
rect 14375 4775 14402 4792
rect 14375 4758 14380 4775
rect 14397 4758 14402 4775
rect 14375 4741 14402 4758
rect 14375 4724 14380 4741
rect 14397 4724 14402 4741
rect 14375 4707 14402 4724
rect 14375 4690 14380 4707
rect 14397 4690 14402 4707
rect 14375 4673 14402 4690
rect 14375 4656 14380 4673
rect 14397 4656 14402 4673
rect 14375 4639 14402 4656
rect 14375 4622 14380 4639
rect 14397 4622 14402 4639
rect 14375 4614 14402 4622
rect 14419 4809 14477 4817
rect 14419 4792 14424 4809
rect 14441 4792 14477 4809
rect 14419 4775 14477 4792
rect 14419 4758 14424 4775
rect 14441 4758 14477 4775
rect 14419 4741 14477 4758
rect 14419 4724 14424 4741
rect 14441 4724 14477 4741
rect 14419 4707 14477 4724
rect 14419 4690 14424 4707
rect 14441 4690 14477 4707
rect 14419 4673 14477 4690
rect 14419 4656 14424 4673
rect 14441 4656 14477 4673
rect 14419 4639 14477 4656
rect 14419 4622 14424 4639
rect 14441 4622 14477 4639
rect 14419 4614 14477 4622
rect 14250 4537 14283 4545
rect 14250 4520 14258 4537
rect 14275 4520 14283 4537
rect 14250 4512 14283 4520
rect 14300 4527 14327 4614
rect 14349 4589 14382 4597
rect 14349 4572 14357 4589
rect 14374 4581 14382 4589
rect 14450 4581 14477 4614
rect 14374 4572 14477 4581
rect 14349 4564 14477 4572
rect 14395 4535 14428 4543
rect 14395 4527 14403 4535
rect 14300 4518 14403 4527
rect 14420 4518 14428 4535
rect 14300 4510 14428 4518
rect 13916 4499 13949 4507
rect 13916 4482 13924 4499
rect 13941 4482 13949 4499
rect 13916 4474 13949 4482
rect 14250 4483 14283 4491
rect 14250 4466 14258 4483
rect 14275 4466 14283 4483
rect 14250 4458 14283 4466
rect 14300 4441 14327 4510
rect 14450 4441 14477 4564
rect 14911 4809 14969 4817
rect 14911 4792 14947 4809
rect 14964 4792 14969 4809
rect 14911 4775 14969 4792
rect 14911 4758 14947 4775
rect 14964 4758 14969 4775
rect 14911 4741 14969 4758
rect 14911 4724 14947 4741
rect 14964 4724 14969 4741
rect 14911 4707 14969 4724
rect 14911 4690 14947 4707
rect 14964 4690 14969 4707
rect 14911 4673 14969 4690
rect 14911 4656 14947 4673
rect 14964 4656 14969 4673
rect 14911 4639 14969 4656
rect 14911 4622 14947 4639
rect 14964 4622 14969 4639
rect 14911 4614 14969 4622
rect 14986 4809 15013 4832
rect 15597 4832 15601 4851
rect 15620 4832 15624 4851
rect 14986 4792 14991 4809
rect 15008 4792 15013 4809
rect 14986 4775 15013 4792
rect 14986 4758 14991 4775
rect 15008 4758 15013 4775
rect 14986 4741 15013 4758
rect 14986 4724 14991 4741
rect 15008 4724 15013 4741
rect 14986 4707 15013 4724
rect 14986 4690 14991 4707
rect 15008 4690 15013 4707
rect 14986 4673 15013 4690
rect 14986 4656 14991 4673
rect 15008 4656 15013 4673
rect 14986 4639 15013 4656
rect 14986 4622 14991 4639
rect 15008 4622 15013 4639
rect 14986 4614 15013 4622
rect 15030 4809 15088 4817
rect 15030 4792 15035 4809
rect 15052 4792 15088 4809
rect 15030 4775 15088 4792
rect 15030 4758 15035 4775
rect 15052 4758 15088 4775
rect 15030 4741 15088 4758
rect 15030 4724 15035 4741
rect 15052 4724 15088 4741
rect 15030 4707 15088 4724
rect 15030 4690 15035 4707
rect 15052 4690 15088 4707
rect 15030 4673 15088 4690
rect 15030 4656 15035 4673
rect 15052 4656 15088 4673
rect 15030 4639 15088 4656
rect 15030 4622 15035 4639
rect 15052 4622 15088 4639
rect 15030 4614 15088 4622
rect 14861 4537 14894 4545
rect 14861 4520 14869 4537
rect 14886 4520 14894 4537
rect 14861 4512 14894 4520
rect 14911 4527 14938 4614
rect 14960 4589 14993 4597
rect 14960 4572 14968 4589
rect 14985 4581 14993 4589
rect 15061 4581 15088 4614
rect 14985 4572 15088 4581
rect 14960 4564 15088 4572
rect 15006 4535 15039 4543
rect 15006 4527 15014 4535
rect 14911 4518 15014 4527
rect 15031 4518 15039 4535
rect 14911 4510 15039 4518
rect 14494 4499 14527 4507
rect 14494 4482 14502 4499
rect 14519 4482 14527 4499
rect 14494 4474 14527 4482
rect 14861 4483 14894 4491
rect 14861 4466 14869 4483
rect 14886 4466 14894 4483
rect 14861 4458 14894 4466
rect 14911 4441 14938 4510
rect 15061 4441 15088 4564
rect 15522 4809 15580 4817
rect 15522 4792 15558 4809
rect 15575 4792 15580 4809
rect 15522 4775 15580 4792
rect 15522 4758 15558 4775
rect 15575 4758 15580 4775
rect 15522 4741 15580 4758
rect 15522 4724 15558 4741
rect 15575 4724 15580 4741
rect 15522 4707 15580 4724
rect 15522 4690 15558 4707
rect 15575 4690 15580 4707
rect 15522 4673 15580 4690
rect 15522 4656 15558 4673
rect 15575 4656 15580 4673
rect 15522 4639 15580 4656
rect 15522 4622 15558 4639
rect 15575 4622 15580 4639
rect 15522 4614 15580 4622
rect 15597 4809 15624 4832
rect 15597 4792 15602 4809
rect 15619 4792 15624 4809
rect 15597 4775 15624 4792
rect 15597 4758 15602 4775
rect 15619 4758 15624 4775
rect 15597 4741 15624 4758
rect 15597 4724 15602 4741
rect 15619 4724 15624 4741
rect 15597 4707 15624 4724
rect 15597 4690 15602 4707
rect 15619 4690 15624 4707
rect 15597 4673 15624 4690
rect 15597 4656 15602 4673
rect 15619 4656 15624 4673
rect 15597 4639 15624 4656
rect 15597 4622 15602 4639
rect 15619 4622 15624 4639
rect 15597 4614 15624 4622
rect 15641 4809 15699 4817
rect 15641 4792 15646 4809
rect 15663 4792 15699 4809
rect 15641 4775 15699 4792
rect 15641 4758 15646 4775
rect 15663 4758 15699 4775
rect 15641 4741 15699 4758
rect 15641 4724 15646 4741
rect 15663 4724 15699 4741
rect 15641 4707 15699 4724
rect 15641 4690 15646 4707
rect 15663 4690 15699 4707
rect 15641 4673 15699 4690
rect 15641 4656 15646 4673
rect 15663 4656 15699 4673
rect 15641 4639 15699 4656
rect 15641 4622 15646 4639
rect 15663 4622 15699 4639
rect 15641 4614 15699 4622
rect 15472 4537 15505 4545
rect 15472 4520 15480 4537
rect 15497 4520 15505 4537
rect 15472 4512 15505 4520
rect 15522 4527 15549 4614
rect 15571 4589 15604 4597
rect 15571 4572 15579 4589
rect 15596 4581 15604 4589
rect 15672 4581 15699 4614
rect 15596 4572 15699 4581
rect 15571 4564 15699 4572
rect 15617 4535 15650 4543
rect 15617 4527 15625 4535
rect 15522 4518 15625 4527
rect 15642 4518 15650 4535
rect 15522 4510 15650 4518
rect 15105 4499 15138 4507
rect 15105 4482 15113 4499
rect 15130 4482 15138 4499
rect 15105 4474 15138 4482
rect 15472 4483 15505 4491
rect 15472 4466 15480 4483
rect 15497 4466 15505 4483
rect 15472 4458 15505 4466
rect 15522 4441 15549 4510
rect 15672 4441 15699 4564
rect 15716 4499 15749 4507
rect 15716 4482 15724 4499
rect 15741 4482 15749 4499
rect 15716 4474 15749 4482
rect 12451 4433 12478 4441
rect 12451 4416 12456 4433
rect 12473 4416 12478 4433
rect 12451 4399 12478 4416
rect 12451 4382 12456 4399
rect 12473 4382 12478 4399
rect 12451 4365 12478 4382
rect 12451 4348 12456 4365
rect 12473 4348 12478 4365
rect 12451 4340 12478 4348
rect 12500 4433 12558 4441
rect 12500 4416 12536 4433
rect 12553 4416 12558 4433
rect 12500 4399 12558 4416
rect 12500 4382 12536 4399
rect 12553 4382 12558 4399
rect 12500 4365 12558 4382
rect 12500 4348 12536 4365
rect 12553 4348 12558 4365
rect 12500 4340 12558 4348
rect 12575 4433 12602 4441
rect 12575 4416 12580 4433
rect 12597 4416 12602 4433
rect 12575 4399 12602 4416
rect 12575 4382 12580 4399
rect 12597 4382 12602 4399
rect 12575 4365 12602 4382
rect 12575 4348 12580 4365
rect 12597 4348 12602 4365
rect 12575 4325 12602 4348
rect 12619 4433 12677 4441
rect 12619 4416 12624 4433
rect 12641 4416 12677 4433
rect 12619 4399 12677 4416
rect 12619 4382 12624 4399
rect 12641 4382 12677 4399
rect 12619 4365 12677 4382
rect 12619 4348 12624 4365
rect 12641 4348 12677 4365
rect 12619 4340 12677 4348
rect 12699 4433 12726 4441
rect 12699 4416 12704 4433
rect 12721 4416 12726 4433
rect 12699 4399 12726 4416
rect 12699 4382 12704 4399
rect 12721 4382 12726 4399
rect 12699 4365 12726 4382
rect 12699 4348 12704 4365
rect 12721 4348 12726 4365
rect 12699 4340 12726 4348
rect 13062 4433 13089 4441
rect 13062 4416 13067 4433
rect 13084 4416 13089 4433
rect 13062 4399 13089 4416
rect 13062 4382 13067 4399
rect 13084 4382 13089 4399
rect 13062 4365 13089 4382
rect 13062 4348 13067 4365
rect 13084 4348 13089 4365
rect 13062 4340 13089 4348
rect 13111 4433 13169 4441
rect 13111 4416 13147 4433
rect 13164 4416 13169 4433
rect 13111 4399 13169 4416
rect 13111 4382 13147 4399
rect 13164 4382 13169 4399
rect 13111 4365 13169 4382
rect 13111 4348 13147 4365
rect 13164 4348 13169 4365
rect 13111 4340 13169 4348
rect 13186 4433 13213 4441
rect 13186 4416 13191 4433
rect 13208 4416 13213 4433
rect 13186 4399 13213 4416
rect 13186 4382 13191 4399
rect 13208 4382 13213 4399
rect 13186 4365 13213 4382
rect 13186 4348 13191 4365
rect 13208 4348 13213 4365
rect 12575 4306 12579 4325
rect 12598 4306 12602 4325
rect 13186 4325 13213 4348
rect 13230 4433 13288 4441
rect 13230 4416 13235 4433
rect 13252 4416 13288 4433
rect 13230 4399 13288 4416
rect 13230 4382 13235 4399
rect 13252 4382 13288 4399
rect 13230 4365 13288 4382
rect 13230 4348 13235 4365
rect 13252 4348 13288 4365
rect 13230 4340 13288 4348
rect 13310 4433 13337 4441
rect 13310 4416 13315 4433
rect 13332 4416 13337 4433
rect 13310 4399 13337 4416
rect 13310 4382 13315 4399
rect 13332 4382 13337 4399
rect 13310 4365 13337 4382
rect 13310 4348 13315 4365
rect 13332 4348 13337 4365
rect 13310 4340 13337 4348
rect 13673 4433 13700 4441
rect 13673 4416 13678 4433
rect 13695 4416 13700 4433
rect 13673 4399 13700 4416
rect 13673 4382 13678 4399
rect 13695 4382 13700 4399
rect 13673 4365 13700 4382
rect 13673 4348 13678 4365
rect 13695 4348 13700 4365
rect 13673 4340 13700 4348
rect 13722 4433 13780 4441
rect 13722 4416 13758 4433
rect 13775 4416 13780 4433
rect 13722 4399 13780 4416
rect 13722 4382 13758 4399
rect 13775 4382 13780 4399
rect 13722 4365 13780 4382
rect 13722 4348 13758 4365
rect 13775 4348 13780 4365
rect 13722 4340 13780 4348
rect 13797 4433 13824 4441
rect 13797 4416 13802 4433
rect 13819 4416 13824 4433
rect 13797 4399 13824 4416
rect 13797 4382 13802 4399
rect 13819 4382 13824 4399
rect 13797 4365 13824 4382
rect 13797 4348 13802 4365
rect 13819 4348 13824 4365
rect 13186 4306 13190 4325
rect 13209 4306 13213 4325
rect 13797 4325 13824 4348
rect 13841 4433 13899 4441
rect 13841 4416 13846 4433
rect 13863 4416 13899 4433
rect 13841 4399 13899 4416
rect 13841 4382 13846 4399
rect 13863 4382 13899 4399
rect 13841 4365 13899 4382
rect 13841 4348 13846 4365
rect 13863 4348 13899 4365
rect 13841 4340 13899 4348
rect 13921 4433 13948 4441
rect 13921 4416 13926 4433
rect 13943 4416 13948 4433
rect 13921 4399 13948 4416
rect 13921 4382 13926 4399
rect 13943 4382 13948 4399
rect 13921 4365 13948 4382
rect 13921 4348 13926 4365
rect 13943 4348 13948 4365
rect 13921 4340 13948 4348
rect 14251 4433 14278 4441
rect 14251 4416 14256 4433
rect 14273 4416 14278 4433
rect 14251 4399 14278 4416
rect 14251 4382 14256 4399
rect 14273 4382 14278 4399
rect 14251 4365 14278 4382
rect 14251 4348 14256 4365
rect 14273 4348 14278 4365
rect 14251 4340 14278 4348
rect 14300 4433 14358 4441
rect 14300 4416 14336 4433
rect 14353 4416 14358 4433
rect 14300 4399 14358 4416
rect 14300 4382 14336 4399
rect 14353 4382 14358 4399
rect 14300 4365 14358 4382
rect 14300 4348 14336 4365
rect 14353 4348 14358 4365
rect 14300 4340 14358 4348
rect 14375 4433 14402 4441
rect 14375 4416 14380 4433
rect 14397 4416 14402 4433
rect 14375 4399 14402 4416
rect 14375 4382 14380 4399
rect 14397 4382 14402 4399
rect 14375 4365 14402 4382
rect 14375 4348 14380 4365
rect 14397 4348 14402 4365
rect 13797 4306 13801 4325
rect 13820 4306 13824 4325
rect 14375 4325 14402 4348
rect 14419 4433 14477 4441
rect 14419 4416 14424 4433
rect 14441 4416 14477 4433
rect 14419 4399 14477 4416
rect 14419 4382 14424 4399
rect 14441 4382 14477 4399
rect 14419 4365 14477 4382
rect 14419 4348 14424 4365
rect 14441 4348 14477 4365
rect 14419 4340 14477 4348
rect 14499 4433 14526 4441
rect 14499 4416 14504 4433
rect 14521 4416 14526 4433
rect 14499 4399 14526 4416
rect 14499 4382 14504 4399
rect 14521 4382 14526 4399
rect 14499 4365 14526 4382
rect 14499 4348 14504 4365
rect 14521 4348 14526 4365
rect 14499 4340 14526 4348
rect 14862 4433 14889 4441
rect 14862 4416 14867 4433
rect 14884 4416 14889 4433
rect 14862 4399 14889 4416
rect 14862 4382 14867 4399
rect 14884 4382 14889 4399
rect 14862 4365 14889 4382
rect 14862 4348 14867 4365
rect 14884 4348 14889 4365
rect 14862 4340 14889 4348
rect 14911 4433 14969 4441
rect 14911 4416 14947 4433
rect 14964 4416 14969 4433
rect 14911 4399 14969 4416
rect 14911 4382 14947 4399
rect 14964 4382 14969 4399
rect 14911 4365 14969 4382
rect 14911 4348 14947 4365
rect 14964 4348 14969 4365
rect 14911 4340 14969 4348
rect 14986 4433 15013 4441
rect 14986 4416 14991 4433
rect 15008 4416 15013 4433
rect 14986 4399 15013 4416
rect 14986 4382 14991 4399
rect 15008 4382 15013 4399
rect 14986 4365 15013 4382
rect 14986 4348 14991 4365
rect 15008 4348 15013 4365
rect 14375 4306 14379 4325
rect 14398 4306 14402 4325
rect 14986 4325 15013 4348
rect 15030 4433 15088 4441
rect 15030 4416 15035 4433
rect 15052 4416 15088 4433
rect 15030 4399 15088 4416
rect 15030 4382 15035 4399
rect 15052 4382 15088 4399
rect 15030 4365 15088 4382
rect 15030 4348 15035 4365
rect 15052 4348 15088 4365
rect 15030 4340 15088 4348
rect 15110 4433 15137 4441
rect 15110 4416 15115 4433
rect 15132 4416 15137 4433
rect 15110 4399 15137 4416
rect 15110 4382 15115 4399
rect 15132 4382 15137 4399
rect 15110 4365 15137 4382
rect 15110 4348 15115 4365
rect 15132 4348 15137 4365
rect 15110 4340 15137 4348
rect 15473 4433 15500 4441
rect 15473 4416 15478 4433
rect 15495 4416 15500 4433
rect 15473 4399 15500 4416
rect 15473 4382 15478 4399
rect 15495 4382 15500 4399
rect 15473 4365 15500 4382
rect 15473 4348 15478 4365
rect 15495 4348 15500 4365
rect 15473 4340 15500 4348
rect 15522 4433 15580 4441
rect 15522 4416 15558 4433
rect 15575 4416 15580 4433
rect 15522 4399 15580 4416
rect 15522 4382 15558 4399
rect 15575 4382 15580 4399
rect 15522 4365 15580 4382
rect 15522 4348 15558 4365
rect 15575 4348 15580 4365
rect 15522 4340 15580 4348
rect 15597 4433 15624 4441
rect 15597 4416 15602 4433
rect 15619 4416 15624 4433
rect 15597 4399 15624 4416
rect 15597 4382 15602 4399
rect 15619 4382 15624 4399
rect 15597 4365 15624 4382
rect 15597 4348 15602 4365
rect 15619 4348 15624 4365
rect 14986 4306 14990 4325
rect 15009 4306 15013 4325
rect 15597 4325 15624 4348
rect 15641 4433 15699 4441
rect 15641 4416 15646 4433
rect 15663 4416 15699 4433
rect 15641 4399 15699 4416
rect 15641 4382 15646 4399
rect 15663 4382 15699 4399
rect 15641 4365 15699 4382
rect 15641 4348 15646 4365
rect 15663 4348 15699 4365
rect 15641 4340 15699 4348
rect 15721 4433 15748 4441
rect 15721 4416 15726 4433
rect 15743 4416 15748 4433
rect 15721 4399 15748 4416
rect 15721 4382 15726 4399
rect 15743 4382 15748 4399
rect 15721 4365 15748 4382
rect 15721 4348 15726 4365
rect 15743 4348 15748 4365
rect 15721 4340 15748 4348
rect 15597 4306 15601 4325
rect 15620 4306 15624 4325
<< viali >>
rect 13190 8062 13209 8081
rect 13801 8062 13820 8081
rect 13069 7750 13086 7767
rect 13168 7802 13185 7819
rect 13214 7748 13231 7765
rect 13069 7696 13086 7713
rect 14379 8062 14398 8081
rect 13680 7750 13697 7767
rect 13779 7802 13796 7819
rect 13825 7748 13842 7765
rect 13313 7712 13330 7729
rect 13680 7696 13697 7713
rect 14990 8062 15009 8081
rect 14258 7750 14275 7767
rect 14357 7802 14374 7819
rect 14403 7748 14420 7765
rect 13924 7712 13941 7729
rect 14258 7696 14275 7713
rect 15601 8062 15620 8081
rect 14869 7750 14886 7767
rect 14968 7802 14985 7819
rect 15014 7748 15031 7765
rect 14502 7712 14519 7729
rect 14869 7696 14886 7713
rect 15480 7750 15497 7767
rect 15579 7802 15596 7819
rect 15625 7748 15642 7765
rect 15113 7712 15130 7729
rect 15480 7696 15497 7713
rect 15724 7712 15741 7729
rect 13190 7536 13209 7555
rect 13801 7536 13820 7555
rect 14379 7536 14398 7555
rect 14990 7536 15009 7555
rect 15601 7536 15620 7555
rect 12579 7412 12598 7431
rect 13190 7412 13209 7431
rect 12458 7100 12475 7117
rect 12557 7152 12574 7169
rect 12603 7098 12620 7115
rect 12458 7046 12475 7063
rect 13801 7412 13820 7431
rect 13069 7100 13086 7117
rect 13168 7152 13185 7169
rect 13214 7098 13231 7115
rect 12702 7062 12719 7079
rect 13069 7046 13086 7063
rect 14379 7412 14398 7431
rect 13680 7100 13697 7117
rect 13779 7152 13796 7169
rect 13825 7098 13842 7115
rect 13313 7062 13330 7079
rect 13680 7046 13697 7063
rect 14990 7412 15009 7431
rect 14258 7100 14275 7117
rect 14357 7152 14374 7169
rect 14403 7098 14420 7115
rect 13924 7062 13941 7079
rect 14258 7046 14275 7063
rect 15601 7412 15620 7431
rect 14869 7100 14886 7117
rect 14968 7152 14985 7169
rect 15014 7098 15031 7115
rect 14502 7062 14519 7079
rect 14869 7046 14886 7063
rect 15480 7100 15497 7117
rect 15579 7152 15596 7169
rect 15625 7098 15642 7115
rect 15113 7062 15130 7079
rect 15480 7046 15497 7063
rect 15724 7062 15741 7079
rect 12579 6886 12598 6905
rect 13190 6886 13209 6905
rect 13801 6886 13820 6905
rect 14379 6886 14398 6905
rect 14990 6886 15009 6905
rect 15601 6886 15620 6905
rect 12579 6772 12598 6791
rect 13190 6772 13209 6791
rect 12458 6460 12475 6477
rect 12557 6512 12574 6529
rect 12603 6458 12620 6475
rect 12458 6406 12475 6423
rect 13801 6772 13820 6791
rect 13069 6460 13086 6477
rect 13168 6512 13185 6529
rect 13214 6458 13231 6475
rect 12702 6422 12719 6439
rect 13069 6406 13086 6423
rect 14379 6772 14398 6791
rect 13680 6460 13697 6477
rect 13779 6512 13796 6529
rect 13825 6458 13842 6475
rect 13313 6422 13330 6439
rect 13680 6406 13697 6423
rect 14990 6772 15009 6791
rect 14258 6460 14275 6477
rect 14357 6512 14374 6529
rect 14403 6458 14420 6475
rect 13924 6422 13941 6439
rect 14258 6406 14275 6423
rect 15601 6772 15620 6791
rect 14869 6460 14886 6477
rect 14968 6512 14985 6529
rect 15014 6458 15031 6475
rect 14502 6422 14519 6439
rect 14869 6406 14886 6423
rect 15480 6460 15497 6477
rect 15579 6512 15596 6529
rect 15625 6458 15642 6475
rect 15113 6422 15130 6439
rect 15480 6406 15497 6423
rect 15724 6422 15741 6439
rect 12579 6246 12598 6265
rect 13190 6246 13209 6265
rect 13801 6246 13820 6265
rect 14379 6246 14398 6265
rect 14990 6246 15009 6265
rect 15601 6246 15620 6265
rect 12579 6122 12598 6141
rect 13190 6122 13209 6141
rect 12458 5810 12475 5827
rect 12557 5862 12574 5879
rect 12603 5808 12620 5825
rect 12458 5756 12475 5773
rect 13801 6122 13820 6141
rect 13069 5810 13086 5827
rect 13168 5862 13185 5879
rect 13214 5808 13231 5825
rect 12702 5772 12719 5789
rect 13069 5756 13086 5773
rect 14379 6122 14398 6141
rect 13680 5810 13697 5827
rect 13779 5862 13796 5879
rect 13825 5808 13842 5825
rect 13313 5772 13330 5789
rect 13680 5756 13697 5773
rect 14990 6122 15009 6141
rect 14258 5810 14275 5827
rect 14357 5862 14374 5879
rect 14403 5808 14420 5825
rect 13924 5772 13941 5789
rect 14258 5756 14275 5773
rect 15601 6122 15620 6141
rect 14869 5810 14886 5827
rect 14968 5862 14985 5879
rect 15014 5808 15031 5825
rect 14502 5772 14519 5789
rect 14869 5756 14886 5773
rect 15480 5810 15497 5827
rect 15579 5862 15596 5879
rect 15625 5808 15642 5825
rect 15113 5772 15130 5789
rect 15480 5756 15497 5773
rect 15724 5772 15741 5789
rect 12579 5596 12598 5615
rect 13190 5596 13209 5615
rect 13801 5596 13820 5615
rect 14379 5596 14398 5615
rect 14990 5596 15009 5615
rect 15601 5596 15620 5615
rect 12579 5472 12598 5491
rect 13190 5472 13209 5491
rect 12458 5160 12475 5177
rect 12557 5212 12574 5229
rect 12603 5158 12620 5175
rect 12458 5106 12475 5123
rect 13801 5472 13820 5491
rect 13069 5160 13086 5177
rect 13168 5212 13185 5229
rect 13214 5158 13231 5175
rect 12702 5122 12719 5139
rect 13069 5106 13086 5123
rect 14379 5472 14398 5491
rect 13680 5160 13697 5177
rect 13779 5212 13796 5229
rect 13825 5158 13842 5175
rect 13313 5122 13330 5139
rect 13680 5106 13697 5123
rect 14990 5472 15009 5491
rect 14258 5160 14275 5177
rect 14357 5212 14374 5229
rect 14403 5158 14420 5175
rect 13924 5122 13941 5139
rect 14258 5106 14275 5123
rect 15601 5472 15620 5491
rect 14869 5160 14886 5177
rect 14968 5212 14985 5229
rect 15014 5158 15031 5175
rect 14502 5122 14519 5139
rect 14869 5106 14886 5123
rect 15480 5160 15497 5177
rect 15579 5212 15596 5229
rect 15625 5158 15642 5175
rect 15113 5122 15130 5139
rect 15480 5106 15497 5123
rect 15724 5122 15741 5139
rect 12579 4946 12598 4965
rect 13190 4946 13209 4965
rect 13801 4946 13820 4965
rect 14379 4946 14398 4965
rect 14990 4946 15009 4965
rect 15601 4946 15620 4965
rect 12579 4832 12598 4851
rect 13190 4832 13209 4851
rect 12458 4520 12475 4537
rect 12557 4572 12574 4589
rect 12603 4518 12620 4535
rect 12458 4466 12475 4483
rect 13801 4832 13820 4851
rect 13069 4520 13086 4537
rect 13168 4572 13185 4589
rect 13214 4518 13231 4535
rect 12702 4482 12719 4499
rect 13069 4466 13086 4483
rect 14379 4832 14398 4851
rect 13680 4520 13697 4537
rect 13779 4572 13796 4589
rect 13825 4518 13842 4535
rect 13313 4482 13330 4499
rect 13680 4466 13697 4483
rect 14990 4832 15009 4851
rect 14258 4520 14275 4537
rect 14357 4572 14374 4589
rect 14403 4518 14420 4535
rect 13924 4482 13941 4499
rect 14258 4466 14275 4483
rect 15601 4832 15620 4851
rect 14869 4520 14886 4537
rect 14968 4572 14985 4589
rect 15014 4518 15031 4535
rect 14502 4482 14519 4499
rect 14869 4466 14886 4483
rect 15480 4520 15497 4537
rect 15579 4572 15596 4589
rect 15625 4518 15642 4535
rect 15113 4482 15130 4499
rect 15480 4466 15497 4483
rect 15724 4482 15741 4499
rect 12579 4306 12598 4325
rect 13190 4306 13209 4325
rect 13801 4306 13820 4325
rect 14379 4306 14398 4325
rect 14990 4306 15009 4325
rect 15601 4306 15620 4325
<< metal1 >>
rect 12280 8081 15891 8096
rect 12280 8062 13190 8081
rect 13209 8062 13801 8081
rect 13820 8062 14379 8081
rect 14398 8062 14990 8081
rect 15009 8062 15601 8081
rect 15620 8062 15891 8081
rect 12280 8047 15891 8062
rect 12518 7824 12582 7827
rect 12518 7797 12521 7824
rect 12548 7797 12582 7824
rect 12518 7794 12582 7797
rect 13160 7819 13193 7827
rect 13160 7802 13168 7819
rect 13185 7802 13193 7819
rect 13160 7794 13193 7802
rect 13771 7819 13804 7827
rect 13771 7802 13779 7819
rect 13796 7802 13804 7819
rect 13771 7794 13804 7802
rect 14318 7824 14382 7827
rect 14318 7797 14321 7824
rect 14348 7819 14382 7824
rect 14348 7802 14357 7819
rect 14374 7802 14382 7819
rect 14348 7797 14382 7802
rect 14318 7794 14382 7797
rect 14960 7819 14993 7827
rect 14960 7802 14968 7819
rect 14985 7802 14993 7819
rect 14960 7794 14993 7802
rect 15571 7819 15604 7827
rect 15571 7802 15579 7819
rect 15596 7802 15604 7819
rect 15571 7794 15604 7802
rect 12302 7771 12483 7775
rect 12302 7745 12305 7771
rect 12331 7745 12483 7771
rect 12302 7742 12483 7745
rect 12595 7770 12661 7773
rect 12595 7743 12631 7770
rect 12658 7743 12661 7770
rect 12595 7740 12661 7743
rect 12913 7771 13094 7775
rect 12913 7745 12916 7771
rect 12942 7767 13094 7771
rect 12942 7750 13069 7767
rect 13086 7750 13094 7767
rect 12942 7745 13094 7750
rect 12913 7742 13094 7745
rect 13206 7765 13239 7773
rect 13206 7748 13214 7765
rect 13231 7748 13239 7765
rect 13206 7740 13239 7748
rect 13524 7771 13705 7775
rect 13524 7745 13527 7771
rect 13553 7767 13705 7771
rect 13553 7750 13680 7767
rect 13697 7750 13705 7767
rect 13553 7745 13705 7750
rect 13524 7742 13705 7745
rect 13817 7765 13850 7773
rect 13817 7748 13825 7765
rect 13842 7748 13850 7765
rect 13817 7740 13850 7748
rect 14102 7771 14283 7775
rect 14102 7745 14105 7771
rect 14131 7767 14283 7771
rect 14131 7750 14258 7767
rect 14275 7750 14283 7767
rect 14131 7745 14283 7750
rect 14102 7742 14283 7745
rect 14395 7770 14461 7773
rect 14395 7765 14431 7770
rect 14395 7748 14403 7765
rect 14420 7748 14431 7765
rect 14395 7743 14431 7748
rect 14458 7743 14461 7770
rect 14395 7740 14461 7743
rect 14713 7771 14894 7775
rect 14713 7745 14716 7771
rect 14742 7767 14894 7771
rect 14742 7750 14869 7767
rect 14886 7750 14894 7767
rect 14742 7745 14894 7750
rect 14713 7742 14894 7745
rect 15006 7765 15039 7773
rect 15006 7748 15014 7765
rect 15031 7748 15039 7765
rect 15006 7740 15039 7748
rect 15324 7771 15505 7775
rect 15324 7745 15327 7771
rect 15353 7767 15505 7771
rect 15353 7750 15480 7767
rect 15497 7750 15505 7767
rect 15353 7745 15505 7750
rect 15324 7742 15505 7745
rect 15617 7765 15650 7773
rect 15617 7748 15625 7765
rect 15642 7748 15650 7765
rect 15617 7740 15650 7748
rect 12694 7733 12805 7737
rect 12402 7717 12483 7721
rect 12402 7691 12405 7717
rect 12431 7691 12483 7717
rect 12694 7707 12775 7733
rect 12801 7707 12805 7733
rect 13305 7733 13416 7737
rect 13305 7729 13386 7733
rect 12694 7704 12805 7707
rect 13013 7717 13094 7721
rect 12402 7688 12483 7691
rect 13013 7691 13016 7717
rect 13042 7713 13094 7717
rect 13042 7696 13069 7713
rect 13086 7696 13094 7713
rect 13305 7712 13313 7729
rect 13330 7712 13386 7729
rect 13305 7707 13386 7712
rect 13412 7707 13416 7733
rect 13916 7733 14027 7737
rect 13916 7729 13997 7733
rect 13305 7704 13416 7707
rect 13624 7717 13705 7721
rect 13042 7691 13094 7696
rect 13013 7688 13094 7691
rect 13624 7691 13627 7717
rect 13653 7713 13705 7717
rect 13653 7696 13680 7713
rect 13697 7696 13705 7713
rect 13916 7712 13924 7729
rect 13941 7712 13997 7729
rect 13916 7707 13997 7712
rect 14023 7707 14027 7733
rect 14494 7733 14605 7737
rect 14494 7729 14575 7733
rect 13916 7704 14027 7707
rect 14202 7717 14283 7721
rect 13653 7691 13705 7696
rect 13624 7688 13705 7691
rect 14202 7691 14205 7717
rect 14231 7713 14283 7717
rect 14231 7696 14258 7713
rect 14275 7696 14283 7713
rect 14494 7712 14502 7729
rect 14519 7712 14575 7729
rect 14494 7707 14575 7712
rect 14601 7707 14605 7733
rect 15105 7733 15216 7737
rect 15105 7729 15186 7733
rect 14494 7704 14605 7707
rect 14813 7717 14894 7721
rect 14231 7691 14283 7696
rect 14202 7688 14283 7691
rect 14813 7691 14816 7717
rect 14842 7713 14894 7717
rect 14842 7696 14869 7713
rect 14886 7696 14894 7713
rect 15105 7712 15113 7729
rect 15130 7712 15186 7729
rect 15105 7707 15186 7712
rect 15212 7707 15216 7733
rect 15716 7733 15827 7737
rect 15716 7729 15797 7733
rect 15105 7704 15216 7707
rect 15424 7717 15505 7721
rect 14842 7691 14894 7696
rect 14813 7688 14894 7691
rect 15424 7691 15427 7717
rect 15453 7713 15505 7717
rect 15453 7696 15480 7713
rect 15497 7696 15505 7713
rect 15716 7712 15724 7729
rect 15741 7712 15797 7729
rect 15716 7707 15797 7712
rect 15823 7707 15827 7733
rect 15716 7704 15827 7707
rect 15453 7691 15505 7696
rect 15424 7688 15505 7691
rect 12247 7555 15891 7570
rect 12247 7536 13190 7555
rect 13209 7536 13801 7555
rect 13820 7536 14379 7555
rect 14398 7536 14990 7555
rect 15009 7536 15601 7555
rect 15620 7536 15891 7555
rect 12247 7521 15891 7536
rect 12261 7431 15891 7446
rect 12261 7412 12579 7431
rect 12598 7412 13190 7431
rect 13209 7412 13801 7431
rect 13820 7412 14379 7431
rect 14398 7412 14990 7431
rect 15009 7412 15601 7431
rect 15620 7412 15891 7431
rect 12261 7397 15891 7412
rect 12516 7174 12582 7177
rect 12516 7147 12519 7174
rect 12546 7169 12582 7174
rect 12546 7152 12557 7169
rect 12574 7152 12582 7169
rect 12546 7147 12582 7152
rect 12516 7144 12582 7147
rect 13127 7173 13193 7177
rect 13127 7146 13133 7173
rect 13160 7169 13193 7173
rect 13160 7152 13168 7169
rect 13185 7152 13193 7169
rect 13160 7146 13193 7152
rect 13127 7144 13193 7146
rect 13738 7173 13804 7177
rect 13738 7146 13743 7173
rect 13770 7169 13804 7173
rect 13770 7152 13779 7169
rect 13796 7152 13804 7169
rect 13770 7146 13804 7152
rect 13738 7144 13804 7146
rect 14316 7174 14382 7177
rect 14316 7147 14319 7174
rect 14346 7169 14382 7174
rect 14346 7152 14357 7169
rect 14374 7152 14382 7169
rect 14346 7147 14382 7152
rect 14316 7144 14382 7147
rect 14927 7173 14993 7177
rect 14927 7146 14933 7173
rect 14960 7169 14993 7173
rect 14960 7152 14968 7169
rect 14985 7152 14993 7169
rect 14960 7146 14993 7152
rect 14927 7144 14993 7146
rect 15538 7173 15604 7177
rect 15538 7146 15543 7173
rect 15570 7169 15604 7173
rect 15570 7152 15579 7169
rect 15596 7152 15604 7169
rect 15570 7146 15604 7152
rect 15538 7144 15604 7146
rect 12302 7121 12483 7125
rect 12302 7095 12305 7121
rect 12331 7117 12483 7121
rect 12331 7100 12458 7117
rect 12475 7100 12483 7117
rect 12331 7095 12483 7100
rect 12302 7092 12483 7095
rect 12595 7120 12661 7123
rect 12595 7115 12631 7120
rect 12595 7098 12603 7115
rect 12620 7098 12631 7115
rect 12595 7093 12631 7098
rect 12658 7093 12661 7120
rect 12595 7090 12661 7093
rect 12913 7121 13094 7125
rect 12913 7095 12916 7121
rect 12942 7117 13094 7121
rect 12942 7100 13069 7117
rect 13086 7100 13094 7117
rect 12942 7095 13094 7100
rect 12913 7092 13094 7095
rect 13206 7120 13266 7123
rect 13206 7115 13239 7120
rect 13206 7098 13214 7115
rect 13231 7098 13239 7115
rect 13206 7093 13239 7098
rect 13206 7090 13266 7093
rect 13524 7121 13705 7125
rect 13524 7095 13527 7121
rect 13553 7117 13705 7121
rect 13553 7100 13680 7117
rect 13697 7100 13705 7117
rect 13553 7095 13705 7100
rect 13524 7092 13705 7095
rect 13817 7120 13882 7123
rect 13817 7115 13851 7120
rect 13817 7098 13825 7115
rect 13842 7098 13851 7115
rect 13817 7093 13851 7098
rect 13878 7093 13882 7120
rect 13817 7090 13882 7093
rect 14102 7121 14283 7125
rect 14102 7095 14105 7121
rect 14131 7117 14283 7121
rect 14131 7100 14258 7117
rect 14275 7100 14283 7117
rect 14131 7095 14283 7100
rect 14102 7092 14283 7095
rect 14395 7120 14461 7123
rect 14395 7115 14431 7120
rect 14395 7098 14403 7115
rect 14420 7098 14431 7115
rect 14395 7093 14431 7098
rect 14458 7093 14461 7120
rect 14395 7090 14461 7093
rect 14713 7121 14894 7125
rect 14713 7095 14716 7121
rect 14742 7117 14894 7121
rect 14742 7100 14869 7117
rect 14886 7100 14894 7117
rect 14742 7095 14894 7100
rect 14713 7092 14894 7095
rect 15006 7120 15066 7123
rect 15006 7115 15039 7120
rect 15006 7098 15014 7115
rect 15031 7098 15039 7115
rect 15006 7093 15039 7098
rect 15006 7090 15066 7093
rect 15324 7121 15505 7125
rect 15324 7095 15327 7121
rect 15353 7117 15505 7121
rect 15353 7100 15480 7117
rect 15497 7100 15505 7117
rect 15353 7095 15505 7100
rect 15324 7092 15505 7095
rect 15617 7120 15682 7123
rect 15617 7115 15651 7120
rect 15617 7098 15625 7115
rect 15642 7098 15651 7115
rect 15617 7093 15651 7098
rect 15678 7093 15682 7120
rect 15617 7090 15682 7093
rect 13234 7089 13266 7090
rect 15034 7089 15066 7090
rect 12694 7083 12805 7087
rect 12694 7079 12775 7083
rect 12402 7067 12483 7071
rect 12402 7041 12405 7067
rect 12431 7063 12483 7067
rect 12431 7046 12458 7063
rect 12475 7046 12483 7063
rect 12694 7062 12702 7079
rect 12719 7062 12775 7079
rect 12694 7057 12775 7062
rect 12801 7057 12805 7083
rect 13305 7083 13416 7087
rect 13305 7079 13386 7083
rect 12694 7054 12805 7057
rect 13013 7067 13094 7071
rect 12431 7041 12483 7046
rect 12402 7038 12483 7041
rect 13013 7041 13016 7067
rect 13042 7063 13094 7067
rect 13042 7046 13069 7063
rect 13086 7046 13094 7063
rect 13305 7062 13313 7079
rect 13330 7062 13386 7079
rect 13305 7057 13386 7062
rect 13412 7057 13416 7083
rect 13916 7083 14027 7087
rect 13916 7079 13997 7083
rect 13305 7054 13416 7057
rect 13624 7067 13705 7071
rect 13042 7041 13094 7046
rect 13013 7038 13094 7041
rect 13624 7041 13627 7067
rect 13653 7063 13705 7067
rect 13653 7046 13680 7063
rect 13697 7046 13705 7063
rect 13916 7062 13924 7079
rect 13941 7062 13997 7079
rect 13916 7057 13997 7062
rect 14023 7057 14027 7083
rect 14494 7083 14605 7087
rect 14494 7079 14575 7083
rect 13916 7054 14027 7057
rect 14202 7067 14283 7071
rect 13653 7041 13705 7046
rect 13624 7038 13705 7041
rect 14202 7041 14205 7067
rect 14231 7063 14283 7067
rect 14231 7046 14258 7063
rect 14275 7046 14283 7063
rect 14494 7062 14502 7079
rect 14519 7062 14575 7079
rect 14494 7057 14575 7062
rect 14601 7057 14605 7083
rect 15105 7083 15216 7087
rect 15105 7079 15186 7083
rect 14494 7054 14605 7057
rect 14813 7067 14894 7071
rect 14231 7041 14283 7046
rect 14202 7038 14283 7041
rect 14813 7041 14816 7067
rect 14842 7063 14894 7067
rect 14842 7046 14869 7063
rect 14886 7046 14894 7063
rect 15105 7062 15113 7079
rect 15130 7062 15186 7079
rect 15105 7057 15186 7062
rect 15212 7057 15216 7083
rect 15716 7083 15827 7087
rect 15716 7079 15797 7083
rect 15105 7054 15216 7057
rect 15424 7067 15505 7071
rect 14842 7041 14894 7046
rect 14813 7038 14894 7041
rect 15424 7041 15427 7067
rect 15453 7063 15505 7067
rect 15453 7046 15480 7063
rect 15497 7046 15505 7063
rect 15716 7062 15724 7079
rect 15741 7062 15797 7079
rect 15716 7057 15797 7062
rect 15823 7057 15827 7083
rect 15716 7054 15827 7057
rect 15453 7041 15505 7046
rect 15424 7038 15505 7041
rect 12235 6905 15891 6920
rect 12235 6886 12579 6905
rect 12598 6886 13190 6905
rect 13209 6886 13801 6905
rect 13820 6886 14379 6905
rect 14398 6886 14990 6905
rect 15009 6886 15601 6905
rect 15620 6886 15891 6905
rect 12235 6871 15891 6886
rect 12253 6791 15891 6806
rect 12253 6772 12579 6791
rect 12598 6772 13190 6791
rect 13209 6772 13801 6791
rect 13820 6772 14379 6791
rect 14398 6772 14990 6791
rect 15009 6772 15601 6791
rect 15620 6772 15891 6791
rect 12253 6757 15891 6772
rect 12516 6534 12582 6537
rect 12516 6507 12519 6534
rect 12546 6529 12582 6534
rect 12546 6512 12557 6529
rect 12574 6512 12582 6529
rect 12546 6507 12582 6512
rect 12516 6504 12582 6507
rect 13128 6534 13193 6537
rect 13128 6507 13133 6534
rect 13160 6529 13193 6534
rect 13160 6512 13168 6529
rect 13185 6512 13193 6529
rect 13160 6507 13193 6512
rect 13128 6504 13193 6507
rect 13739 6534 13804 6537
rect 13739 6507 13744 6534
rect 13771 6529 13804 6534
rect 13771 6512 13779 6529
rect 13796 6512 13804 6529
rect 13771 6507 13804 6512
rect 13739 6504 13804 6507
rect 14316 6534 14382 6537
rect 14316 6507 14319 6534
rect 14346 6529 14382 6534
rect 14346 6512 14357 6529
rect 14374 6512 14382 6529
rect 14346 6507 14382 6512
rect 14316 6504 14382 6507
rect 14928 6534 14993 6537
rect 14928 6507 14933 6534
rect 14960 6529 14993 6534
rect 14960 6512 14968 6529
rect 14985 6512 14993 6529
rect 14960 6507 14993 6512
rect 14928 6504 14993 6507
rect 15539 6534 15604 6537
rect 15539 6507 15544 6534
rect 15571 6529 15604 6534
rect 15571 6512 15579 6529
rect 15596 6512 15604 6529
rect 15571 6507 15604 6512
rect 15539 6504 15604 6507
rect 12302 6481 12483 6485
rect 12302 6455 12305 6481
rect 12331 6477 12483 6481
rect 12331 6460 12458 6477
rect 12475 6460 12483 6477
rect 12331 6455 12483 6460
rect 12302 6452 12483 6455
rect 12595 6480 12661 6483
rect 12595 6475 12631 6480
rect 12595 6458 12603 6475
rect 12620 6458 12631 6475
rect 12595 6453 12631 6458
rect 12658 6453 12661 6480
rect 12595 6450 12661 6453
rect 12913 6481 13094 6485
rect 12913 6455 12916 6481
rect 12942 6477 13094 6481
rect 12942 6460 13069 6477
rect 13086 6460 13094 6477
rect 12942 6455 13094 6460
rect 12913 6452 13094 6455
rect 13206 6480 13271 6483
rect 13206 6475 13239 6480
rect 13206 6458 13214 6475
rect 13231 6458 13239 6475
rect 13206 6453 13239 6458
rect 13266 6453 13271 6480
rect 13206 6450 13271 6453
rect 13524 6481 13705 6485
rect 13524 6455 13527 6481
rect 13553 6477 13705 6481
rect 13553 6460 13680 6477
rect 13697 6460 13705 6477
rect 13553 6455 13705 6460
rect 13524 6452 13705 6455
rect 13817 6480 13882 6483
rect 13817 6475 13850 6480
rect 13817 6458 13825 6475
rect 13842 6458 13850 6475
rect 13817 6453 13850 6458
rect 13877 6453 13882 6480
rect 13817 6450 13882 6453
rect 14102 6481 14283 6485
rect 14102 6455 14105 6481
rect 14131 6477 14283 6481
rect 14131 6460 14258 6477
rect 14275 6460 14283 6477
rect 14131 6455 14283 6460
rect 14102 6452 14283 6455
rect 14395 6480 14461 6483
rect 14395 6475 14431 6480
rect 14395 6458 14403 6475
rect 14420 6458 14431 6475
rect 14395 6453 14431 6458
rect 14458 6453 14461 6480
rect 14395 6450 14461 6453
rect 14713 6481 14894 6485
rect 14713 6455 14716 6481
rect 14742 6477 14894 6481
rect 14742 6460 14869 6477
rect 14886 6460 14894 6477
rect 14742 6455 14894 6460
rect 14713 6452 14894 6455
rect 15006 6480 15071 6483
rect 15006 6475 15039 6480
rect 15006 6458 15014 6475
rect 15031 6458 15039 6475
rect 15006 6453 15039 6458
rect 15066 6453 15071 6480
rect 15006 6450 15071 6453
rect 15324 6481 15505 6485
rect 15324 6455 15327 6481
rect 15353 6477 15505 6481
rect 15353 6460 15480 6477
rect 15497 6460 15505 6477
rect 15353 6455 15505 6460
rect 15324 6452 15505 6455
rect 15617 6480 15682 6483
rect 15617 6475 15650 6480
rect 15617 6458 15625 6475
rect 15642 6458 15650 6475
rect 15617 6453 15650 6458
rect 15677 6453 15682 6480
rect 15617 6450 15682 6453
rect 12694 6443 12805 6447
rect 12694 6439 12775 6443
rect 12402 6427 12483 6431
rect 12402 6401 12405 6427
rect 12431 6423 12483 6427
rect 12431 6406 12458 6423
rect 12475 6406 12483 6423
rect 12694 6422 12702 6439
rect 12719 6422 12775 6439
rect 12694 6417 12775 6422
rect 12801 6417 12805 6443
rect 13305 6443 13416 6447
rect 13305 6439 13386 6443
rect 12694 6414 12805 6417
rect 13013 6427 13094 6431
rect 12431 6401 12483 6406
rect 12402 6398 12483 6401
rect 13013 6401 13016 6427
rect 13042 6423 13094 6427
rect 13042 6406 13069 6423
rect 13086 6406 13094 6423
rect 13305 6422 13313 6439
rect 13330 6422 13386 6439
rect 13305 6417 13386 6422
rect 13412 6417 13416 6443
rect 13916 6443 14027 6447
rect 13916 6439 13997 6443
rect 13305 6414 13416 6417
rect 13624 6427 13705 6431
rect 13042 6401 13094 6406
rect 13013 6398 13094 6401
rect 13624 6401 13627 6427
rect 13653 6423 13705 6427
rect 13653 6406 13680 6423
rect 13697 6406 13705 6423
rect 13916 6422 13924 6439
rect 13941 6422 13997 6439
rect 13916 6417 13997 6422
rect 14023 6417 14027 6443
rect 14494 6443 14605 6447
rect 14494 6439 14575 6443
rect 13916 6414 14027 6417
rect 14202 6427 14283 6431
rect 13653 6401 13705 6406
rect 13624 6398 13705 6401
rect 14202 6401 14205 6427
rect 14231 6423 14283 6427
rect 14231 6406 14258 6423
rect 14275 6406 14283 6423
rect 14494 6422 14502 6439
rect 14519 6422 14575 6439
rect 14494 6417 14575 6422
rect 14601 6417 14605 6443
rect 15105 6443 15216 6447
rect 15105 6439 15186 6443
rect 14494 6414 14605 6417
rect 14813 6427 14894 6431
rect 14231 6401 14283 6406
rect 14202 6398 14283 6401
rect 14813 6401 14816 6427
rect 14842 6423 14894 6427
rect 14842 6406 14869 6423
rect 14886 6406 14894 6423
rect 15105 6422 15113 6439
rect 15130 6422 15186 6439
rect 15105 6417 15186 6422
rect 15212 6417 15216 6443
rect 15716 6443 15827 6447
rect 15716 6439 15797 6443
rect 15105 6414 15216 6417
rect 15424 6427 15505 6431
rect 14842 6401 14894 6406
rect 14813 6398 14894 6401
rect 15424 6401 15427 6427
rect 15453 6423 15505 6427
rect 15453 6406 15480 6423
rect 15497 6406 15505 6423
rect 15716 6422 15724 6439
rect 15741 6422 15797 6439
rect 15716 6417 15797 6422
rect 15823 6417 15827 6443
rect 15716 6414 15827 6417
rect 15453 6401 15505 6406
rect 15424 6398 15505 6401
rect 12275 6265 15891 6280
rect 12275 6246 12579 6265
rect 12598 6246 13190 6265
rect 13209 6246 13801 6265
rect 13820 6246 14379 6265
rect 14398 6246 14990 6265
rect 15009 6246 15601 6265
rect 15620 6246 15891 6265
rect 12275 6231 15891 6246
rect 12280 6141 15891 6156
rect 12280 6122 12579 6141
rect 12598 6122 13190 6141
rect 13209 6122 13801 6141
rect 13820 6122 14379 6141
rect 14398 6122 14990 6141
rect 15009 6122 15601 6141
rect 15620 6122 15891 6141
rect 12280 6107 15891 6122
rect 12518 5884 12582 5887
rect 12518 5857 12521 5884
rect 12548 5879 12582 5884
rect 12548 5862 12557 5879
rect 12574 5862 12582 5879
rect 12548 5857 12582 5862
rect 12518 5854 12582 5857
rect 13160 5879 13193 5887
rect 13160 5862 13168 5879
rect 13185 5862 13193 5879
rect 13160 5854 13193 5862
rect 13771 5879 13804 5887
rect 13771 5862 13779 5879
rect 13796 5862 13804 5879
rect 13771 5854 13804 5862
rect 14318 5884 14382 5887
rect 14318 5857 14321 5884
rect 14348 5879 14382 5884
rect 14348 5862 14357 5879
rect 14374 5862 14382 5879
rect 14348 5857 14382 5862
rect 14318 5854 14382 5857
rect 14960 5879 14993 5887
rect 14960 5862 14968 5879
rect 14985 5862 14993 5879
rect 14960 5854 14993 5862
rect 15571 5879 15604 5887
rect 15571 5862 15579 5879
rect 15596 5862 15604 5879
rect 15571 5854 15604 5862
rect 12302 5831 12483 5835
rect 12302 5805 12305 5831
rect 12331 5827 12483 5831
rect 12331 5810 12458 5827
rect 12475 5810 12483 5827
rect 12331 5805 12483 5810
rect 12302 5802 12483 5805
rect 12595 5830 12661 5833
rect 12595 5825 12631 5830
rect 12595 5808 12603 5825
rect 12620 5808 12631 5825
rect 12595 5803 12631 5808
rect 12658 5803 12661 5830
rect 12595 5800 12661 5803
rect 12913 5831 13094 5835
rect 12913 5805 12916 5831
rect 12942 5827 13094 5831
rect 12942 5810 13069 5827
rect 13086 5810 13094 5827
rect 12942 5805 13094 5810
rect 12913 5802 13094 5805
rect 13206 5825 13239 5833
rect 13206 5808 13214 5825
rect 13231 5808 13239 5825
rect 13206 5800 13239 5808
rect 13524 5831 13705 5835
rect 13524 5805 13527 5831
rect 13553 5827 13705 5831
rect 13553 5810 13680 5827
rect 13697 5810 13705 5827
rect 13553 5805 13705 5810
rect 13524 5802 13705 5805
rect 13817 5825 13850 5833
rect 13817 5808 13825 5825
rect 13842 5808 13850 5825
rect 13817 5800 13850 5808
rect 14102 5831 14283 5835
rect 14102 5805 14105 5831
rect 14131 5827 14283 5831
rect 14131 5810 14258 5827
rect 14275 5810 14283 5827
rect 14131 5805 14283 5810
rect 14102 5802 14283 5805
rect 14395 5830 14461 5833
rect 14395 5825 14431 5830
rect 14395 5808 14403 5825
rect 14420 5808 14431 5825
rect 14395 5803 14431 5808
rect 14458 5803 14461 5830
rect 14395 5800 14461 5803
rect 14713 5831 14894 5835
rect 14713 5805 14716 5831
rect 14742 5827 14894 5831
rect 14742 5810 14869 5827
rect 14886 5810 14894 5827
rect 14742 5805 14894 5810
rect 14713 5802 14894 5805
rect 15006 5825 15039 5833
rect 15006 5808 15014 5825
rect 15031 5808 15039 5825
rect 15006 5800 15039 5808
rect 15324 5831 15505 5835
rect 15324 5805 15327 5831
rect 15353 5827 15505 5831
rect 15353 5810 15480 5827
rect 15497 5810 15505 5827
rect 15353 5805 15505 5810
rect 15324 5802 15505 5805
rect 15617 5825 15650 5833
rect 15617 5808 15625 5825
rect 15642 5808 15650 5825
rect 15617 5800 15650 5808
rect 12694 5793 12805 5797
rect 12694 5789 12775 5793
rect 12402 5777 12483 5781
rect 12402 5751 12405 5777
rect 12431 5773 12483 5777
rect 12431 5756 12458 5773
rect 12475 5756 12483 5773
rect 12694 5772 12702 5789
rect 12719 5772 12775 5789
rect 12694 5767 12775 5772
rect 12801 5767 12805 5793
rect 13305 5793 13416 5797
rect 13305 5789 13386 5793
rect 12694 5764 12805 5767
rect 13013 5777 13094 5781
rect 12431 5751 12483 5756
rect 12402 5748 12483 5751
rect 13013 5751 13016 5777
rect 13042 5773 13094 5777
rect 13042 5756 13069 5773
rect 13086 5756 13094 5773
rect 13305 5772 13313 5789
rect 13330 5772 13386 5789
rect 13305 5767 13386 5772
rect 13412 5767 13416 5793
rect 13916 5793 14027 5797
rect 13916 5789 13997 5793
rect 13305 5764 13416 5767
rect 13624 5777 13705 5781
rect 13042 5751 13094 5756
rect 13013 5748 13094 5751
rect 13624 5751 13627 5777
rect 13653 5773 13705 5777
rect 13653 5756 13680 5773
rect 13697 5756 13705 5773
rect 13916 5772 13924 5789
rect 13941 5772 13997 5789
rect 13916 5767 13997 5772
rect 14023 5767 14027 5793
rect 14494 5793 14605 5797
rect 14494 5789 14575 5793
rect 13916 5764 14027 5767
rect 14202 5777 14283 5781
rect 13653 5751 13705 5756
rect 13624 5748 13705 5751
rect 14202 5751 14205 5777
rect 14231 5773 14283 5777
rect 14231 5756 14258 5773
rect 14275 5756 14283 5773
rect 14494 5772 14502 5789
rect 14519 5772 14575 5789
rect 14494 5767 14575 5772
rect 14601 5767 14605 5793
rect 15105 5793 15216 5797
rect 15105 5789 15186 5793
rect 14494 5764 14605 5767
rect 14813 5777 14894 5781
rect 14231 5751 14283 5756
rect 14202 5748 14283 5751
rect 14813 5751 14816 5777
rect 14842 5773 14894 5777
rect 14842 5756 14869 5773
rect 14886 5756 14894 5773
rect 15105 5772 15113 5789
rect 15130 5772 15186 5789
rect 15105 5767 15186 5772
rect 15212 5767 15216 5793
rect 15716 5793 15827 5797
rect 15716 5789 15797 5793
rect 15105 5764 15216 5767
rect 15424 5777 15505 5781
rect 14842 5751 14894 5756
rect 14813 5748 14894 5751
rect 15424 5751 15427 5777
rect 15453 5773 15505 5777
rect 15453 5756 15480 5773
rect 15497 5756 15505 5773
rect 15716 5772 15724 5789
rect 15741 5772 15797 5789
rect 15716 5767 15797 5772
rect 15823 5767 15827 5793
rect 15716 5764 15827 5767
rect 15453 5751 15505 5756
rect 15424 5748 15505 5751
rect 12247 5615 15891 5630
rect 12247 5596 12579 5615
rect 12598 5596 13190 5615
rect 13209 5596 13801 5615
rect 13820 5596 14379 5615
rect 14398 5596 14990 5615
rect 15009 5596 15601 5615
rect 15620 5596 15891 5615
rect 12247 5581 15891 5596
rect 12261 5491 15891 5506
rect 12261 5472 12579 5491
rect 12598 5472 13190 5491
rect 13209 5472 13801 5491
rect 13820 5472 14379 5491
rect 14398 5472 14990 5491
rect 15009 5472 15601 5491
rect 15620 5472 15891 5491
rect 12261 5457 15891 5472
rect 12516 5234 12582 5237
rect 12516 5207 12519 5234
rect 12546 5229 12582 5234
rect 12546 5212 12557 5229
rect 12574 5212 12582 5229
rect 12546 5207 12582 5212
rect 12516 5204 12582 5207
rect 13127 5233 13193 5237
rect 13127 5206 13133 5233
rect 13160 5229 13193 5233
rect 13160 5212 13168 5229
rect 13185 5212 13193 5229
rect 13160 5206 13193 5212
rect 13127 5204 13193 5206
rect 13738 5233 13804 5237
rect 13738 5206 13743 5233
rect 13770 5229 13804 5233
rect 13770 5212 13779 5229
rect 13796 5212 13804 5229
rect 13770 5206 13804 5212
rect 13738 5204 13804 5206
rect 14316 5234 14382 5237
rect 14316 5207 14319 5234
rect 14346 5229 14382 5234
rect 14346 5212 14357 5229
rect 14374 5212 14382 5229
rect 14346 5207 14382 5212
rect 14316 5204 14382 5207
rect 14927 5233 14993 5237
rect 14927 5206 14933 5233
rect 14960 5229 14993 5233
rect 14960 5212 14968 5229
rect 14985 5212 14993 5229
rect 14960 5206 14993 5212
rect 14927 5204 14993 5206
rect 15538 5233 15604 5237
rect 15538 5206 15543 5233
rect 15570 5229 15604 5233
rect 15570 5212 15579 5229
rect 15596 5212 15604 5229
rect 15570 5206 15604 5212
rect 15538 5204 15604 5206
rect 12302 5181 12483 5185
rect 12302 5155 12305 5181
rect 12331 5177 12483 5181
rect 12331 5160 12458 5177
rect 12475 5160 12483 5177
rect 12331 5155 12483 5160
rect 12302 5152 12483 5155
rect 12595 5180 12661 5183
rect 12595 5175 12631 5180
rect 12595 5158 12603 5175
rect 12620 5158 12631 5175
rect 12595 5153 12631 5158
rect 12658 5153 12661 5180
rect 12595 5150 12661 5153
rect 12913 5181 13094 5185
rect 12913 5155 12916 5181
rect 12942 5177 13094 5181
rect 12942 5160 13069 5177
rect 13086 5160 13094 5177
rect 12942 5155 13094 5160
rect 12913 5152 13094 5155
rect 13206 5180 13266 5183
rect 13206 5175 13239 5180
rect 13206 5158 13214 5175
rect 13231 5158 13239 5175
rect 13206 5153 13239 5158
rect 13206 5150 13266 5153
rect 13524 5181 13705 5185
rect 13524 5155 13527 5181
rect 13553 5177 13705 5181
rect 13553 5160 13680 5177
rect 13697 5160 13705 5177
rect 13553 5155 13705 5160
rect 13524 5152 13705 5155
rect 13817 5180 13882 5183
rect 13817 5175 13851 5180
rect 13817 5158 13825 5175
rect 13842 5158 13851 5175
rect 13817 5153 13851 5158
rect 13878 5153 13882 5180
rect 13817 5150 13882 5153
rect 14102 5181 14283 5185
rect 14102 5155 14105 5181
rect 14131 5177 14283 5181
rect 14131 5160 14258 5177
rect 14275 5160 14283 5177
rect 14131 5155 14283 5160
rect 14102 5152 14283 5155
rect 14395 5180 14461 5183
rect 14395 5175 14431 5180
rect 14395 5158 14403 5175
rect 14420 5158 14431 5175
rect 14395 5153 14431 5158
rect 14458 5153 14461 5180
rect 14395 5150 14461 5153
rect 14713 5181 14894 5185
rect 14713 5155 14716 5181
rect 14742 5177 14894 5181
rect 14742 5160 14869 5177
rect 14886 5160 14894 5177
rect 14742 5155 14894 5160
rect 14713 5152 14894 5155
rect 15006 5180 15066 5183
rect 15006 5175 15039 5180
rect 15006 5158 15014 5175
rect 15031 5158 15039 5175
rect 15006 5153 15039 5158
rect 15006 5150 15066 5153
rect 15324 5181 15505 5185
rect 15324 5155 15327 5181
rect 15353 5177 15505 5181
rect 15353 5160 15480 5177
rect 15497 5160 15505 5177
rect 15353 5155 15505 5160
rect 15324 5152 15505 5155
rect 15617 5180 15682 5183
rect 15617 5175 15651 5180
rect 15617 5158 15625 5175
rect 15642 5158 15651 5175
rect 15617 5153 15651 5158
rect 15678 5153 15682 5180
rect 15617 5150 15682 5153
rect 13234 5149 13266 5150
rect 15034 5149 15066 5150
rect 12694 5143 12805 5147
rect 12694 5139 12775 5143
rect 12402 5127 12483 5131
rect 12402 5101 12405 5127
rect 12431 5123 12483 5127
rect 12431 5106 12458 5123
rect 12475 5106 12483 5123
rect 12694 5122 12702 5139
rect 12719 5122 12775 5139
rect 12694 5117 12775 5122
rect 12801 5117 12805 5143
rect 13305 5143 13416 5147
rect 13305 5139 13386 5143
rect 12694 5114 12805 5117
rect 13013 5127 13094 5131
rect 12431 5101 12483 5106
rect 12402 5098 12483 5101
rect 13013 5101 13016 5127
rect 13042 5123 13094 5127
rect 13042 5106 13069 5123
rect 13086 5106 13094 5123
rect 13305 5122 13313 5139
rect 13330 5122 13386 5139
rect 13305 5117 13386 5122
rect 13412 5117 13416 5143
rect 13916 5143 14027 5147
rect 13916 5139 13997 5143
rect 13305 5114 13416 5117
rect 13624 5127 13705 5131
rect 13042 5101 13094 5106
rect 13013 5098 13094 5101
rect 13624 5101 13627 5127
rect 13653 5123 13705 5127
rect 13653 5106 13680 5123
rect 13697 5106 13705 5123
rect 13916 5122 13924 5139
rect 13941 5122 13997 5139
rect 13916 5117 13997 5122
rect 14023 5117 14027 5143
rect 14494 5143 14605 5147
rect 14494 5139 14575 5143
rect 13916 5114 14027 5117
rect 14202 5127 14283 5131
rect 13653 5101 13705 5106
rect 13624 5098 13705 5101
rect 14202 5101 14205 5127
rect 14231 5123 14283 5127
rect 14231 5106 14258 5123
rect 14275 5106 14283 5123
rect 14494 5122 14502 5139
rect 14519 5122 14575 5139
rect 14494 5117 14575 5122
rect 14601 5117 14605 5143
rect 15105 5143 15216 5147
rect 15105 5139 15186 5143
rect 14494 5114 14605 5117
rect 14813 5127 14894 5131
rect 14231 5101 14283 5106
rect 14202 5098 14283 5101
rect 14813 5101 14816 5127
rect 14842 5123 14894 5127
rect 14842 5106 14869 5123
rect 14886 5106 14894 5123
rect 15105 5122 15113 5139
rect 15130 5122 15186 5139
rect 15105 5117 15186 5122
rect 15212 5117 15216 5143
rect 15716 5143 15827 5147
rect 15716 5139 15797 5143
rect 15105 5114 15216 5117
rect 15424 5127 15505 5131
rect 14842 5101 14894 5106
rect 14813 5098 14894 5101
rect 15424 5101 15427 5127
rect 15453 5123 15505 5127
rect 15453 5106 15480 5123
rect 15497 5106 15505 5123
rect 15716 5122 15724 5139
rect 15741 5122 15797 5139
rect 15716 5117 15797 5122
rect 15823 5117 15827 5143
rect 15716 5114 15827 5117
rect 15453 5101 15505 5106
rect 15424 5098 15505 5101
rect 12235 4965 15891 4980
rect 12235 4946 12579 4965
rect 12598 4946 13190 4965
rect 13209 4946 13801 4965
rect 13820 4946 14379 4965
rect 14398 4946 14990 4965
rect 15009 4946 15601 4965
rect 15620 4946 15891 4965
rect 12235 4931 15891 4946
rect 12253 4851 15891 4866
rect 12253 4832 12579 4851
rect 12598 4832 13190 4851
rect 13209 4832 13801 4851
rect 13820 4832 14379 4851
rect 14398 4832 14990 4851
rect 15009 4832 15601 4851
rect 15620 4832 15891 4851
rect 12253 4817 15891 4832
rect 12516 4594 12582 4597
rect 12516 4567 12519 4594
rect 12546 4589 12582 4594
rect 12546 4572 12557 4589
rect 12574 4572 12582 4589
rect 12546 4567 12582 4572
rect 12516 4564 12582 4567
rect 13128 4594 13193 4597
rect 13128 4567 13133 4594
rect 13160 4589 13193 4594
rect 13160 4572 13168 4589
rect 13185 4572 13193 4589
rect 13160 4567 13193 4572
rect 13128 4564 13193 4567
rect 13739 4594 13804 4597
rect 13739 4567 13744 4594
rect 13771 4589 13804 4594
rect 13771 4572 13779 4589
rect 13796 4572 13804 4589
rect 13771 4567 13804 4572
rect 13739 4564 13804 4567
rect 14316 4594 14382 4597
rect 14316 4567 14319 4594
rect 14346 4589 14382 4594
rect 14346 4572 14357 4589
rect 14374 4572 14382 4589
rect 14346 4567 14382 4572
rect 14316 4564 14382 4567
rect 14928 4594 14993 4597
rect 14928 4567 14933 4594
rect 14960 4589 14993 4594
rect 14960 4572 14968 4589
rect 14985 4572 14993 4589
rect 14960 4567 14993 4572
rect 14928 4564 14993 4567
rect 15539 4594 15604 4597
rect 15539 4567 15544 4594
rect 15571 4589 15604 4594
rect 15571 4572 15579 4589
rect 15596 4572 15604 4589
rect 15571 4567 15604 4572
rect 15539 4564 15604 4567
rect 12302 4541 12483 4545
rect 12302 4515 12305 4541
rect 12331 4537 12483 4541
rect 12331 4520 12458 4537
rect 12475 4520 12483 4537
rect 12331 4515 12483 4520
rect 12302 4512 12483 4515
rect 12595 4540 12661 4543
rect 12595 4535 12631 4540
rect 12595 4518 12603 4535
rect 12620 4518 12631 4535
rect 12595 4513 12631 4518
rect 12658 4513 12661 4540
rect 12595 4510 12661 4513
rect 12913 4541 13094 4545
rect 12913 4515 12916 4541
rect 12942 4537 13094 4541
rect 12942 4520 13069 4537
rect 13086 4520 13094 4537
rect 12942 4515 13094 4520
rect 12913 4512 13094 4515
rect 13206 4540 13271 4543
rect 13206 4535 13239 4540
rect 13206 4518 13214 4535
rect 13231 4518 13239 4535
rect 13206 4513 13239 4518
rect 13266 4513 13271 4540
rect 13206 4510 13271 4513
rect 13524 4541 13705 4545
rect 13524 4515 13527 4541
rect 13553 4537 13705 4541
rect 13553 4520 13680 4537
rect 13697 4520 13705 4537
rect 13553 4515 13705 4520
rect 13524 4512 13705 4515
rect 13817 4540 13882 4543
rect 13817 4535 13850 4540
rect 13817 4518 13825 4535
rect 13842 4518 13850 4535
rect 13817 4513 13850 4518
rect 13877 4513 13882 4540
rect 13817 4510 13882 4513
rect 14102 4541 14283 4545
rect 14102 4515 14105 4541
rect 14131 4537 14283 4541
rect 14131 4520 14258 4537
rect 14275 4520 14283 4537
rect 14131 4515 14283 4520
rect 14102 4512 14283 4515
rect 14395 4540 14461 4543
rect 14395 4535 14431 4540
rect 14395 4518 14403 4535
rect 14420 4518 14431 4535
rect 14395 4513 14431 4518
rect 14458 4513 14461 4540
rect 14395 4510 14461 4513
rect 14713 4541 14894 4545
rect 14713 4515 14716 4541
rect 14742 4537 14894 4541
rect 14742 4520 14869 4537
rect 14886 4520 14894 4537
rect 14742 4515 14894 4520
rect 14713 4512 14894 4515
rect 15006 4540 15071 4543
rect 15006 4535 15039 4540
rect 15006 4518 15014 4535
rect 15031 4518 15039 4535
rect 15006 4513 15039 4518
rect 15066 4513 15071 4540
rect 15006 4510 15071 4513
rect 15324 4541 15505 4545
rect 15324 4515 15327 4541
rect 15353 4537 15505 4541
rect 15353 4520 15480 4537
rect 15497 4520 15505 4537
rect 15353 4515 15505 4520
rect 15324 4512 15505 4515
rect 15617 4540 15682 4543
rect 15617 4535 15650 4540
rect 15617 4518 15625 4535
rect 15642 4518 15650 4535
rect 15617 4513 15650 4518
rect 15677 4513 15682 4540
rect 15617 4510 15682 4513
rect 12694 4503 12805 4507
rect 12694 4499 12775 4503
rect 12402 4487 12483 4491
rect 12402 4461 12405 4487
rect 12431 4483 12483 4487
rect 12431 4466 12458 4483
rect 12475 4466 12483 4483
rect 12694 4482 12702 4499
rect 12719 4482 12775 4499
rect 12694 4477 12775 4482
rect 12801 4477 12805 4503
rect 13305 4503 13416 4507
rect 13305 4499 13386 4503
rect 12694 4474 12805 4477
rect 13013 4487 13094 4491
rect 12431 4461 12483 4466
rect 12402 4458 12483 4461
rect 13013 4461 13016 4487
rect 13042 4483 13094 4487
rect 13042 4466 13069 4483
rect 13086 4466 13094 4483
rect 13305 4482 13313 4499
rect 13330 4482 13386 4499
rect 13305 4477 13386 4482
rect 13412 4477 13416 4503
rect 13916 4503 14027 4507
rect 13916 4499 13997 4503
rect 13305 4474 13416 4477
rect 13624 4487 13705 4491
rect 13042 4461 13094 4466
rect 13013 4458 13094 4461
rect 13624 4461 13627 4487
rect 13653 4483 13705 4487
rect 13653 4466 13680 4483
rect 13697 4466 13705 4483
rect 13916 4482 13924 4499
rect 13941 4482 13997 4499
rect 13916 4477 13997 4482
rect 14023 4477 14027 4503
rect 14494 4503 14605 4507
rect 14494 4499 14575 4503
rect 13916 4474 14027 4477
rect 14202 4487 14283 4491
rect 13653 4461 13705 4466
rect 13624 4458 13705 4461
rect 14202 4461 14205 4487
rect 14231 4483 14283 4487
rect 14231 4466 14258 4483
rect 14275 4466 14283 4483
rect 14494 4482 14502 4499
rect 14519 4482 14575 4499
rect 14494 4477 14575 4482
rect 14601 4477 14605 4503
rect 15105 4503 15216 4507
rect 15105 4499 15186 4503
rect 14494 4474 14605 4477
rect 14813 4487 14894 4491
rect 14231 4461 14283 4466
rect 14202 4458 14283 4461
rect 14813 4461 14816 4487
rect 14842 4483 14894 4487
rect 14842 4466 14869 4483
rect 14886 4466 14894 4483
rect 15105 4482 15113 4499
rect 15130 4482 15186 4499
rect 15105 4477 15186 4482
rect 15212 4477 15216 4503
rect 15716 4503 15827 4507
rect 15716 4499 15797 4503
rect 15105 4474 15216 4477
rect 15424 4487 15505 4491
rect 14842 4461 14894 4466
rect 14813 4458 14894 4461
rect 15424 4461 15427 4487
rect 15453 4483 15505 4487
rect 15453 4466 15480 4483
rect 15497 4466 15505 4483
rect 15716 4482 15724 4499
rect 15741 4482 15797 4499
rect 15716 4477 15797 4482
rect 15823 4477 15827 4503
rect 15716 4474 15827 4477
rect 15453 4461 15505 4466
rect 15424 4458 15505 4461
rect 12275 4325 15891 4340
rect 12275 4306 12579 4325
rect 12598 4306 13190 4325
rect 13209 4306 13801 4325
rect 13820 4306 14379 4325
rect 14398 4306 14990 4325
rect 15009 4306 15601 4325
rect 15620 4306 15891 4325
rect 12275 4291 15891 4306
rect 975 1218 14336 1266
rect 975 1156 1025 1218
rect 600 1155 1025 1156
rect 251 1154 1025 1155
rect 100 1145 1025 1154
rect 100 1113 154 1145
rect 186 1113 1025 1145
rect 100 1105 1025 1113
rect 100 1104 400 1105
rect 13249 890 14137 915
rect 13249 850 13274 890
rect 13314 850 14137 890
rect 13249 825 14137 850
rect 14267 890 15271 915
rect 14267 850 15206 890
rect 15246 850 15271 890
rect 14267 825 15271 850
rect 400 633 14335 683
<< via1 >>
rect 12521 7797 12548 7824
rect 14321 7797 14348 7824
rect 12305 7745 12331 7771
rect 12631 7743 12658 7770
rect 12916 7745 12942 7771
rect 13527 7745 13553 7771
rect 14105 7745 14131 7771
rect 14431 7743 14458 7770
rect 14716 7745 14742 7771
rect 15327 7745 15353 7771
rect 12405 7691 12431 7717
rect 12775 7707 12801 7733
rect 13016 7691 13042 7717
rect 13386 7707 13412 7733
rect 13627 7691 13653 7717
rect 13997 7707 14023 7733
rect 14205 7691 14231 7717
rect 14575 7707 14601 7733
rect 14816 7691 14842 7717
rect 15186 7707 15212 7733
rect 15427 7691 15453 7717
rect 15797 7707 15823 7733
rect 12519 7147 12546 7174
rect 13133 7146 13160 7173
rect 13743 7146 13770 7173
rect 14319 7147 14346 7174
rect 14933 7146 14960 7173
rect 15543 7146 15570 7173
rect 12305 7095 12331 7121
rect 12631 7093 12658 7120
rect 12916 7095 12942 7121
rect 13239 7093 13266 7120
rect 13527 7095 13553 7121
rect 13851 7093 13878 7120
rect 14105 7095 14131 7121
rect 14431 7093 14458 7120
rect 14716 7095 14742 7121
rect 15039 7093 15066 7120
rect 15327 7095 15353 7121
rect 15651 7093 15678 7120
rect 12405 7041 12431 7067
rect 12775 7057 12801 7083
rect 13016 7041 13042 7067
rect 13386 7057 13412 7083
rect 13627 7041 13653 7067
rect 13997 7057 14023 7083
rect 14205 7041 14231 7067
rect 14575 7057 14601 7083
rect 14816 7041 14842 7067
rect 15186 7057 15212 7083
rect 15427 7041 15453 7067
rect 15797 7057 15823 7083
rect 12519 6507 12546 6534
rect 13133 6507 13160 6534
rect 13744 6507 13771 6534
rect 14319 6507 14346 6534
rect 14933 6507 14960 6534
rect 15544 6507 15571 6534
rect 12305 6455 12331 6481
rect 12631 6453 12658 6480
rect 12916 6455 12942 6481
rect 13239 6453 13266 6480
rect 13527 6455 13553 6481
rect 13850 6453 13877 6480
rect 14105 6455 14131 6481
rect 14431 6453 14458 6480
rect 14716 6455 14742 6481
rect 15039 6453 15066 6480
rect 15327 6455 15353 6481
rect 15650 6453 15677 6480
rect 12405 6401 12431 6427
rect 12775 6417 12801 6443
rect 13016 6401 13042 6427
rect 13386 6417 13412 6443
rect 13627 6401 13653 6427
rect 13997 6417 14023 6443
rect 14205 6401 14231 6427
rect 14575 6417 14601 6443
rect 14816 6401 14842 6427
rect 15186 6417 15212 6443
rect 15427 6401 15453 6427
rect 15797 6417 15823 6443
rect 12521 5857 12548 5884
rect 14321 5857 14348 5884
rect 12305 5805 12331 5831
rect 12631 5803 12658 5830
rect 12916 5805 12942 5831
rect 13527 5805 13553 5831
rect 14105 5805 14131 5831
rect 14431 5803 14458 5830
rect 14716 5805 14742 5831
rect 15327 5805 15353 5831
rect 12405 5751 12431 5777
rect 12775 5767 12801 5793
rect 13016 5751 13042 5777
rect 13386 5767 13412 5793
rect 13627 5751 13653 5777
rect 13997 5767 14023 5793
rect 14205 5751 14231 5777
rect 14575 5767 14601 5793
rect 14816 5751 14842 5777
rect 15186 5767 15212 5793
rect 15427 5751 15453 5777
rect 15797 5767 15823 5793
rect 12519 5207 12546 5234
rect 13133 5206 13160 5233
rect 13743 5206 13770 5233
rect 14319 5207 14346 5234
rect 14933 5206 14960 5233
rect 15543 5206 15570 5233
rect 12305 5155 12331 5181
rect 12631 5153 12658 5180
rect 12916 5155 12942 5181
rect 13239 5153 13266 5180
rect 13527 5155 13553 5181
rect 13851 5153 13878 5180
rect 14105 5155 14131 5181
rect 14431 5153 14458 5180
rect 14716 5155 14742 5181
rect 15039 5153 15066 5180
rect 15327 5155 15353 5181
rect 15651 5153 15678 5180
rect 12405 5101 12431 5127
rect 12775 5117 12801 5143
rect 13016 5101 13042 5127
rect 13386 5117 13412 5143
rect 13627 5101 13653 5127
rect 13997 5117 14023 5143
rect 14205 5101 14231 5127
rect 14575 5117 14601 5143
rect 14816 5101 14842 5127
rect 15186 5117 15212 5143
rect 15427 5101 15453 5127
rect 15797 5117 15823 5143
rect 12519 4567 12546 4594
rect 13133 4567 13160 4594
rect 13744 4567 13771 4594
rect 14319 4567 14346 4594
rect 14933 4567 14960 4594
rect 15544 4567 15571 4594
rect 12305 4515 12331 4541
rect 12631 4513 12658 4540
rect 12916 4515 12942 4541
rect 13239 4513 13266 4540
rect 13527 4515 13553 4541
rect 13850 4513 13877 4540
rect 14105 4515 14131 4541
rect 14431 4513 14458 4540
rect 14716 4515 14742 4541
rect 15039 4513 15066 4540
rect 15327 4515 15353 4541
rect 15650 4513 15677 4540
rect 12405 4461 12431 4487
rect 12775 4477 12801 4503
rect 13016 4461 13042 4487
rect 13386 4477 13412 4503
rect 13627 4461 13653 4487
rect 13997 4477 14023 4503
rect 14205 4461 14231 4487
rect 14575 4477 14601 4503
rect 14816 4461 14842 4487
rect 15186 4477 15212 4503
rect 15427 4461 15453 4487
rect 15797 4477 15823 4503
rect 154 1113 186 1145
rect 13274 850 13314 890
rect 15206 850 15246 890
<< metal2 >>
rect 12302 7771 12335 8136
rect 12302 7745 12305 7771
rect 12331 7745 12335 7771
rect 12302 7121 12335 7745
rect 12302 7095 12305 7121
rect 12331 7095 12335 7121
rect 12302 6481 12335 7095
rect 12302 6455 12305 6481
rect 12331 6455 12335 6481
rect 12302 5831 12335 6455
rect 12302 5805 12305 5831
rect 12331 5805 12335 5831
rect 12302 5181 12335 5805
rect 12302 5155 12305 5181
rect 12331 5155 12335 5181
rect 12302 4541 12335 5155
rect 12302 4515 12305 4541
rect 12331 4515 12335 4541
rect 12302 4247 12335 4515
rect 12402 7717 12435 8136
rect 12402 7691 12405 7717
rect 12431 7691 12435 7717
rect 12402 7067 12435 7691
rect 12518 7824 12553 8136
rect 12518 7797 12521 7824
rect 12548 7797 12553 7824
rect 12518 7177 12553 7797
rect 12516 7174 12553 7177
rect 12516 7147 12519 7174
rect 12546 7147 12553 7174
rect 12516 7144 12553 7147
rect 12402 7041 12405 7067
rect 12431 7041 12435 7067
rect 12402 6427 12435 7041
rect 12518 6537 12553 7144
rect 12402 6401 12405 6427
rect 12431 6401 12435 6427
rect 12402 5777 12435 6401
rect 12516 6534 12553 6537
rect 12516 6507 12519 6534
rect 12546 6507 12553 6534
rect 12516 6188 12553 6507
rect 12402 5751 12405 5777
rect 12431 5751 12435 5777
rect 12402 5127 12435 5751
rect 12518 5884 12553 6188
rect 12518 5857 12521 5884
rect 12548 5857 12553 5884
rect 12518 5237 12553 5857
rect 12516 5234 12553 5237
rect 12516 5207 12519 5234
rect 12546 5207 12553 5234
rect 12516 5204 12553 5207
rect 12402 5101 12405 5127
rect 12431 5101 12435 5127
rect 12402 4487 12435 5101
rect 12518 4597 12553 5204
rect 12402 4461 12405 4487
rect 12431 4461 12435 4487
rect 12402 4247 12435 4461
rect 12516 4594 12553 4597
rect 12516 4567 12519 4594
rect 12546 4567 12553 4594
rect 12516 4248 12553 4567
rect 12624 7770 12661 8136
rect 12624 7743 12631 7770
rect 12658 7743 12661 7770
rect 12624 7120 12661 7743
rect 12624 7093 12631 7120
rect 12658 7093 12661 7120
rect 12624 6480 12661 7093
rect 12624 6453 12631 6480
rect 12658 6453 12661 6480
rect 12624 5830 12661 6453
rect 12624 5803 12631 5830
rect 12658 5803 12661 5830
rect 12624 5180 12661 5803
rect 12624 5153 12631 5180
rect 12658 5153 12661 5180
rect 12624 4540 12661 5153
rect 12624 4513 12631 4540
rect 12658 4513 12661 4540
rect 12624 4245 12661 4513
rect 12772 7733 12805 8136
rect 12772 7707 12775 7733
rect 12801 7707 12805 7733
rect 12772 7083 12805 7707
rect 12772 7057 12775 7083
rect 12801 7057 12805 7083
rect 12772 6443 12805 7057
rect 12772 6417 12775 6443
rect 12801 6417 12805 6443
rect 12772 5793 12805 6417
rect 12772 5767 12775 5793
rect 12801 5767 12805 5793
rect 12772 5143 12805 5767
rect 12772 5117 12775 5143
rect 12801 5117 12805 5143
rect 12772 4503 12805 5117
rect 12772 4477 12775 4503
rect 12801 4477 12805 4503
rect 12772 4247 12805 4477
rect 12913 7771 12946 8136
rect 12913 7745 12916 7771
rect 12942 7745 12946 7771
rect 12913 7121 12946 7745
rect 12913 7095 12916 7121
rect 12942 7095 12946 7121
rect 12913 6481 12946 7095
rect 12913 6455 12916 6481
rect 12942 6455 12946 6481
rect 12913 5831 12946 6455
rect 12913 5805 12916 5831
rect 12942 5805 12946 5831
rect 12913 5181 12946 5805
rect 12913 5155 12916 5181
rect 12942 5155 12946 5181
rect 12913 4541 12946 5155
rect 12913 4515 12916 4541
rect 12942 4515 12946 4541
rect 12913 4247 12946 4515
rect 13013 7717 13046 8136
rect 13013 7691 13016 7717
rect 13042 7691 13046 7717
rect 13013 7067 13046 7691
rect 13013 7041 13016 7067
rect 13042 7041 13046 7067
rect 13013 6427 13046 7041
rect 13013 6401 13016 6427
rect 13042 6401 13046 6427
rect 13013 5777 13046 6401
rect 13013 5751 13016 5777
rect 13042 5751 13046 5777
rect 13013 5127 13046 5751
rect 13013 5101 13016 5127
rect 13042 5101 13046 5127
rect 13013 4487 13046 5101
rect 13013 4461 13016 4487
rect 13042 4461 13046 4487
rect 13013 4247 13046 4461
rect 13127 7173 13164 8136
rect 13127 7146 13133 7173
rect 13160 7146 13164 7173
rect 13127 6534 13164 7146
rect 13127 6507 13133 6534
rect 13160 6507 13164 6534
rect 13127 5233 13164 6507
rect 13127 5206 13133 5233
rect 13160 5206 13164 5233
rect 13127 4594 13164 5206
rect 13127 4567 13133 4594
rect 13160 4567 13164 4594
rect 13127 4250 13164 4567
rect 13235 7120 13272 8136
rect 13235 7093 13239 7120
rect 13266 7093 13272 7120
rect 13235 6480 13272 7093
rect 13235 6453 13239 6480
rect 13266 6453 13272 6480
rect 13235 5180 13272 6453
rect 13235 5153 13239 5180
rect 13266 5153 13272 5180
rect 13235 4540 13272 5153
rect 13235 4513 13239 4540
rect 13266 4513 13272 4540
rect 13235 4253 13272 4513
rect 13383 7733 13416 8136
rect 13383 7707 13386 7733
rect 13412 7707 13416 7733
rect 13383 7083 13416 7707
rect 13383 7057 13386 7083
rect 13412 7057 13416 7083
rect 13383 6443 13416 7057
rect 13383 6417 13386 6443
rect 13412 6417 13416 6443
rect 13383 5793 13416 6417
rect 13383 5767 13386 5793
rect 13412 5767 13416 5793
rect 13383 5143 13416 5767
rect 13383 5117 13386 5143
rect 13412 5117 13416 5143
rect 13383 4503 13416 5117
rect 13383 4477 13386 4503
rect 13412 4477 13416 4503
rect 13383 4247 13416 4477
rect 13524 7771 13557 8136
rect 13524 7745 13527 7771
rect 13553 7745 13557 7771
rect 13524 7121 13557 7745
rect 13524 7095 13527 7121
rect 13553 7095 13557 7121
rect 13524 6481 13557 7095
rect 13524 6455 13527 6481
rect 13553 6455 13557 6481
rect 13524 5831 13557 6455
rect 13524 5805 13527 5831
rect 13553 5805 13557 5831
rect 13524 5181 13557 5805
rect 13524 5155 13527 5181
rect 13553 5155 13557 5181
rect 13524 4541 13557 5155
rect 13524 4515 13527 4541
rect 13553 4515 13557 4541
rect 13524 4247 13557 4515
rect 13624 7717 13657 8136
rect 13624 7691 13627 7717
rect 13653 7691 13657 7717
rect 13624 7067 13657 7691
rect 13624 7041 13627 7067
rect 13653 7041 13657 7067
rect 13624 6427 13657 7041
rect 13624 6401 13627 6427
rect 13653 6401 13657 6427
rect 13624 5777 13657 6401
rect 13624 5751 13627 5777
rect 13653 5751 13657 5777
rect 13624 5127 13657 5751
rect 13624 5101 13627 5127
rect 13653 5101 13657 5127
rect 13624 4487 13657 5101
rect 13624 4461 13627 4487
rect 13653 4461 13657 4487
rect 13624 4247 13657 4461
rect 13738 7173 13775 8136
rect 13738 7146 13743 7173
rect 13770 7146 13775 7173
rect 13738 6534 13775 7146
rect 13738 6507 13744 6534
rect 13771 6507 13775 6534
rect 13738 5233 13775 6507
rect 13738 5206 13743 5233
rect 13770 5206 13775 5233
rect 13738 4594 13775 5206
rect 13738 4567 13744 4594
rect 13771 4567 13775 4594
rect 13738 4251 13775 4567
rect 13846 7120 13883 8136
rect 13846 7093 13851 7120
rect 13878 7093 13883 7120
rect 13846 6480 13883 7093
rect 13846 6453 13850 6480
rect 13877 6453 13883 6480
rect 13846 5180 13883 6453
rect 13846 5153 13851 5180
rect 13878 5153 13883 5180
rect 13846 4540 13883 5153
rect 13846 4513 13850 4540
rect 13877 4513 13883 4540
rect 13846 4252 13883 4513
rect 13994 7733 14027 8136
rect 13994 7707 13997 7733
rect 14023 7707 14027 7733
rect 13994 7083 14027 7707
rect 13994 7057 13997 7083
rect 14023 7057 14027 7083
rect 13994 6443 14027 7057
rect 13994 6417 13997 6443
rect 14023 6417 14027 6443
rect 13994 5793 14027 6417
rect 13994 5767 13997 5793
rect 14023 5767 14027 5793
rect 13994 5143 14027 5767
rect 13994 5117 13997 5143
rect 14023 5117 14027 5143
rect 13994 4503 14027 5117
rect 13994 4477 13997 4503
rect 14023 4477 14027 4503
rect 13994 4247 14027 4477
rect 14102 7771 14135 8136
rect 14102 7745 14105 7771
rect 14131 7745 14135 7771
rect 14102 7121 14135 7745
rect 14102 7095 14105 7121
rect 14131 7095 14135 7121
rect 14102 6481 14135 7095
rect 14102 6455 14105 6481
rect 14131 6455 14135 6481
rect 14102 5831 14135 6455
rect 14102 5805 14105 5831
rect 14131 5805 14135 5831
rect 14102 5181 14135 5805
rect 14102 5155 14105 5181
rect 14131 5155 14135 5181
rect 14102 4541 14135 5155
rect 14102 4515 14105 4541
rect 14131 4515 14135 4541
rect 14102 4247 14135 4515
rect 14202 7717 14235 8136
rect 14202 7691 14205 7717
rect 14231 7691 14235 7717
rect 14202 7067 14235 7691
rect 14318 7824 14353 8136
rect 14318 7797 14321 7824
rect 14348 7797 14353 7824
rect 14318 7177 14353 7797
rect 14316 7174 14353 7177
rect 14316 7147 14319 7174
rect 14346 7147 14353 7174
rect 14316 7144 14353 7147
rect 14202 7041 14205 7067
rect 14231 7041 14235 7067
rect 14202 6427 14235 7041
rect 14318 6537 14353 7144
rect 14202 6401 14205 6427
rect 14231 6401 14235 6427
rect 14202 5777 14235 6401
rect 14316 6534 14353 6537
rect 14316 6507 14319 6534
rect 14346 6507 14353 6534
rect 14316 6188 14353 6507
rect 14202 5751 14205 5777
rect 14231 5751 14235 5777
rect 14202 5127 14235 5751
rect 14318 5884 14353 6188
rect 14318 5857 14321 5884
rect 14348 5857 14353 5884
rect 14318 5237 14353 5857
rect 14316 5234 14353 5237
rect 14316 5207 14319 5234
rect 14346 5207 14353 5234
rect 14316 5204 14353 5207
rect 14202 5101 14205 5127
rect 14231 5101 14235 5127
rect 14202 4487 14235 5101
rect 14318 4597 14353 5204
rect 14202 4461 14205 4487
rect 14231 4461 14235 4487
rect 14202 4247 14235 4461
rect 14316 4594 14353 4597
rect 14316 4567 14319 4594
rect 14346 4567 14353 4594
rect 14316 4248 14353 4567
rect 14424 7770 14461 8136
rect 14424 7743 14431 7770
rect 14458 7743 14461 7770
rect 14424 7120 14461 7743
rect 14424 7093 14431 7120
rect 14458 7093 14461 7120
rect 14424 6480 14461 7093
rect 14424 6453 14431 6480
rect 14458 6453 14461 6480
rect 14424 5830 14461 6453
rect 14424 5803 14431 5830
rect 14458 5803 14461 5830
rect 14424 5180 14461 5803
rect 14424 5153 14431 5180
rect 14458 5153 14461 5180
rect 14424 4540 14461 5153
rect 14424 4513 14431 4540
rect 14458 4513 14461 4540
rect 14424 4245 14461 4513
rect 14572 7733 14605 8136
rect 14572 7707 14575 7733
rect 14601 7707 14605 7733
rect 14572 7083 14605 7707
rect 14572 7057 14575 7083
rect 14601 7057 14605 7083
rect 14572 6443 14605 7057
rect 14572 6417 14575 6443
rect 14601 6417 14605 6443
rect 14572 5793 14605 6417
rect 14572 5767 14575 5793
rect 14601 5767 14605 5793
rect 14572 5143 14605 5767
rect 14572 5117 14575 5143
rect 14601 5117 14605 5143
rect 14572 4503 14605 5117
rect 14572 4477 14575 4503
rect 14601 4477 14605 4503
rect 14572 4247 14605 4477
rect 14713 7771 14746 8136
rect 14713 7745 14716 7771
rect 14742 7745 14746 7771
rect 14713 7121 14746 7745
rect 14713 7095 14716 7121
rect 14742 7095 14746 7121
rect 14713 6481 14746 7095
rect 14713 6455 14716 6481
rect 14742 6455 14746 6481
rect 14713 5831 14746 6455
rect 14713 5805 14716 5831
rect 14742 5805 14746 5831
rect 14713 5181 14746 5805
rect 14713 5155 14716 5181
rect 14742 5155 14746 5181
rect 14713 4541 14746 5155
rect 14713 4515 14716 4541
rect 14742 4515 14746 4541
rect 14713 4247 14746 4515
rect 14813 7717 14846 8136
rect 14813 7691 14816 7717
rect 14842 7691 14846 7717
rect 14813 7067 14846 7691
rect 14813 7041 14816 7067
rect 14842 7041 14846 7067
rect 14813 6427 14846 7041
rect 14813 6401 14816 6427
rect 14842 6401 14846 6427
rect 14813 5777 14846 6401
rect 14813 5751 14816 5777
rect 14842 5751 14846 5777
rect 14813 5127 14846 5751
rect 14813 5101 14816 5127
rect 14842 5101 14846 5127
rect 14813 4487 14846 5101
rect 14813 4461 14816 4487
rect 14842 4461 14846 4487
rect 14813 4247 14846 4461
rect 14927 7173 14964 8136
rect 14927 7146 14933 7173
rect 14960 7146 14964 7173
rect 14927 6534 14964 7146
rect 14927 6507 14933 6534
rect 14960 6507 14964 6534
rect 14927 5233 14964 6507
rect 14927 5206 14933 5233
rect 14960 5206 14964 5233
rect 14927 4594 14964 5206
rect 14927 4567 14933 4594
rect 14960 4567 14964 4594
rect 14927 4250 14964 4567
rect 15035 7120 15072 8136
rect 15035 7093 15039 7120
rect 15066 7093 15072 7120
rect 15035 6480 15072 7093
rect 15035 6453 15039 6480
rect 15066 6453 15072 6480
rect 15035 5180 15072 6453
rect 15035 5153 15039 5180
rect 15066 5153 15072 5180
rect 15035 4540 15072 5153
rect 15035 4513 15039 4540
rect 15066 4513 15072 4540
rect 15035 4253 15072 4513
rect 15183 7733 15216 8136
rect 15183 7707 15186 7733
rect 15212 7707 15216 7733
rect 15183 7083 15216 7707
rect 15183 7057 15186 7083
rect 15212 7057 15216 7083
rect 15183 6443 15216 7057
rect 15183 6417 15186 6443
rect 15212 6417 15216 6443
rect 15183 5793 15216 6417
rect 15183 5767 15186 5793
rect 15212 5767 15216 5793
rect 15183 5143 15216 5767
rect 15183 5117 15186 5143
rect 15212 5117 15216 5143
rect 15183 4503 15216 5117
rect 15183 4477 15186 4503
rect 15212 4477 15216 4503
rect 15183 4247 15216 4477
rect 15324 7771 15357 8136
rect 15324 7745 15327 7771
rect 15353 7745 15357 7771
rect 15324 7121 15357 7745
rect 15324 7095 15327 7121
rect 15353 7095 15357 7121
rect 15324 6481 15357 7095
rect 15324 6455 15327 6481
rect 15353 6455 15357 6481
rect 15324 5831 15357 6455
rect 15324 5805 15327 5831
rect 15353 5805 15357 5831
rect 15324 5181 15357 5805
rect 15324 5155 15327 5181
rect 15353 5155 15357 5181
rect 15324 4541 15357 5155
rect 15324 4515 15327 4541
rect 15353 4515 15357 4541
rect 15324 4247 15357 4515
rect 15424 7717 15457 8136
rect 15424 7691 15427 7717
rect 15453 7691 15457 7717
rect 15424 7067 15457 7691
rect 15424 7041 15427 7067
rect 15453 7041 15457 7067
rect 15424 6427 15457 7041
rect 15424 6401 15427 6427
rect 15453 6401 15457 6427
rect 15424 5777 15457 6401
rect 15424 5751 15427 5777
rect 15453 5751 15457 5777
rect 15424 5127 15457 5751
rect 15424 5101 15427 5127
rect 15453 5101 15457 5127
rect 15424 4487 15457 5101
rect 15424 4461 15427 4487
rect 15453 4461 15457 4487
rect 15424 4247 15457 4461
rect 15538 7173 15575 8136
rect 15538 7146 15543 7173
rect 15570 7146 15575 7173
rect 15538 6534 15575 7146
rect 15538 6507 15544 6534
rect 15571 6507 15575 6534
rect 15538 5233 15575 6507
rect 15538 5206 15543 5233
rect 15570 5206 15575 5233
rect 15538 4594 15575 5206
rect 15538 4567 15544 4594
rect 15571 4567 15575 4594
rect 15538 4251 15575 4567
rect 15646 7120 15683 8136
rect 15646 7093 15651 7120
rect 15678 7093 15683 7120
rect 15646 6480 15683 7093
rect 15646 6453 15650 6480
rect 15677 6453 15683 6480
rect 15646 5180 15683 6453
rect 15646 5153 15651 5180
rect 15678 5153 15683 5180
rect 15646 4540 15683 5153
rect 15646 4513 15650 4540
rect 15677 4513 15683 4540
rect 15646 4252 15683 4513
rect 15794 7733 15827 8136
rect 15794 7707 15797 7733
rect 15823 7707 15827 7733
rect 15794 7083 15827 7707
rect 15794 7057 15797 7083
rect 15823 7057 15827 7083
rect 15794 6443 15827 7057
rect 15794 6417 15797 6443
rect 15823 6417 15827 6443
rect 15794 5793 15827 6417
rect 15794 5767 15797 5793
rect 15823 5767 15827 5793
rect 15794 5143 15827 5767
rect 15794 5117 15797 5143
rect 15823 5117 15827 5143
rect 15794 4503 15827 5117
rect 15794 4477 15797 4503
rect 15823 4477 15827 4503
rect 15794 4247 15827 4477
rect 100 1145 300 1154
rect 100 1113 154 1145
rect 186 1113 300 1145
rect 100 1104 300 1113
rect 13249 890 13339 915
rect 13249 850 13274 890
rect 13314 850 13339 890
rect 13249 825 13339 850
rect 15181 890 15271 915
rect 15181 850 15206 890
rect 15246 850 15271 890
rect 15181 825 15271 850
rect 400 674 600 683
rect 400 642 466 674
rect 498 642 600 674
rect 400 633 600 642
<< via2 >>
rect 154 1113 186 1145
rect 13274 850 13314 890
rect 15206 850 15246 890
rect 466 642 498 674
<< metal3 >>
rect 100 1145 300 1154
rect 100 1113 154 1145
rect 186 1113 300 1145
rect 100 1104 300 1113
rect 13249 890 13339 915
rect 13249 850 13274 890
rect 13314 850 13339 890
rect 13249 825 13339 850
rect 15181 890 15271 915
rect 15181 850 15206 890
rect 15246 850 15271 890
rect 15181 825 15271 850
rect 400 674 600 683
rect 400 642 466 674
rect 498 642 600 674
rect 400 633 600 642
<< via3 >>
rect 154 1113 186 1145
rect 13274 850 13314 890
rect 15206 850 15246 890
rect 466 642 498 674
<< metal4 >>
rect 3067 22476 3097 22576
rect 3343 22476 3373 22576
rect 3619 22476 3649 22576
rect 3895 22476 3925 22576
rect 4171 22476 4201 22576
rect 4447 22476 4477 22576
rect 4723 22476 4753 22576
rect 4999 22476 5029 22576
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 7483 22476 7513 22576
rect 7759 22476 7789 22576
rect 8035 22476 8065 22576
rect 8311 22476 8341 22576
rect 8587 22476 8617 22576
rect 8863 22476 8893 22576
rect 9139 22476 9169 22576
rect 9415 22476 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 100 1145 300 22076
rect 100 1113 154 1145
rect 186 1113 300 1145
rect 100 500 300 1113
rect 400 674 600 22076
rect 400 642 466 674
rect 498 642 600 674
rect 400 500 600 642
rect 13249 890 13339 915
rect 13249 850 13274 890
rect 13314 850 13339 890
rect 1657 0 1747 100
rect 3589 0 3679 100
rect 5521 0 5611 100
rect 7453 0 7543 100
rect 9385 0 9475 100
rect 11317 0 11407 100
rect 13249 0 13339 850
rect 15181 890 15271 915
rect 15181 850 15206 890
rect 15246 850 15271 890
rect 15181 0 15271 850
use latch_sr  latch_sr_0
timestamp 1753205587
transform 1 0 12452 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_1
timestamp 1753205587
transform 1 0 12452 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_2
timestamp 1753205587
transform 1 0 12452 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_3
timestamp 1753205587
transform 1 0 13063 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_4
timestamp 1753205587
transform 1 0 13063 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_5
timestamp 1753205587
transform 1 0 13063 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_6
timestamp 1753205587
transform 1 0 13674 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_7
timestamp 1753205587
transform 1 0 13674 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_8
timestamp 1753205587
transform 1 0 13674 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_9
timestamp 1753205587
transform 1 0 14252 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_10
timestamp 1753205587
transform 1 0 14863 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_11
timestamp 1753205587
transform 1 0 15474 0 1 6280
box -2 -49 275 526
use latch_sr  latch_sr_12
timestamp 1753205587
transform 1 0 14252 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_13
timestamp 1753205587
transform 1 0 14863 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_14
timestamp 1753205587
transform 1 0 15474 0 1 6920
box -2 -49 275 526
use latch_sr  latch_sr_15
timestamp 1753205587
transform 1 0 14252 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_16
timestamp 1753205587
transform 1 0 14863 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_17
timestamp 1753205587
transform 1 0 15474 0 1 7570
box -2 -49 275 526
use latch_sr  latch_sr_18
timestamp 1753205587
transform 1 0 15474 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_19
timestamp 1753205587
transform 1 0 14863 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_20
timestamp 1753205587
transform 1 0 14252 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_21
timestamp 1753205587
transform 1 0 13674 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_22
timestamp 1753205587
transform 1 0 13063 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_23
timestamp 1753205587
transform 1 0 12452 0 1 5630
box -2 -49 275 526
use latch_sr  latch_sr_24
timestamp 1753205587
transform 1 0 15474 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_25
timestamp 1753205587
transform 1 0 14863 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_26
timestamp 1753205587
transform 1 0 14252 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_27
timestamp 1753205587
transform 1 0 13674 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_28
timestamp 1753205587
transform 1 0 13063 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_29
timestamp 1753205587
transform 1 0 12452 0 1 4980
box -2 -49 275 526
use latch_sr  latch_sr_30
timestamp 1753205587
transform 1 0 15474 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_31
timestamp 1753205587
transform 1 0 14863 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_32
timestamp 1753205587
transform 1 0 14252 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_33
timestamp 1753205587
transform 1 0 13674 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_34
timestamp 1753205587
transform 1 0 13063 0 1 4340
box -2 -49 275 526
use latch_sr  latch_sr_35
timestamp 1753205587
transform 1 0 12452 0 1 4340
box -2 -49 275 526
use NOT  NOT_0
timestamp 1750779130
transform 1 0 14171 0 1 657
box -87 -24 160 609
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 15181 0 15271 100 0 FreeSans 480 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 13249 0 13339 100 0 FreeSans 480 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 11317 0 11407 100 0 FreeSans 480 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 9385 0 9475 100 0 FreeSans 480 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 7453 0 7543 100 0 FreeSans 480 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 5521 0 5611 100 0 FreeSans 480 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 3589 0 3679 100 0 FreeSans 480 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 1657 0 1747 100 0 FreeSans 480 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 100 500 300 22076 1 FreeSans 200 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 200 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
