VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOT
  CLASS CORE ;
  FOREIGN NOT ;
  ORIGIN 0.190 0.240 ;
  SIZE 1.790 BY 3.200 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT -0.190 1.080 0.630 1.280 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.426400 ;
    PORT
      LAYER li1 ;
        RECT 0.720 1.490 1.050 2.460 ;
        RECT 0.800 1.280 1.050 1.490 ;
        RECT 0.800 1.080 1.600 1.280 ;
        RECT 0.800 0.890 1.050 1.080 ;
        RECT 0.720 0.260 1.050 0.890 ;
    END
  END Y
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.630 1.380 2.810 ;
        RECT 0.320 1.490 0.550 2.630 ;
      LAYER met1 ;
        RECT -0.190 2.480 1.600 2.960 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.320 0.090 0.550 0.910 ;
        RECT 0.000 -0.090 1.380 0.090 ;
      LAYER met1 ;
        RECT -0.190 -0.240 1.600 0.240 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT -0.190 1.300 1.600 2.910 ;
      LAYER pwell ;
        RECT 0.210 0.890 0.720 1.020 ;
        RECT 0.800 0.890 1.140 1.020 ;
        RECT 0.210 -0.090 1.140 0.890 ;
  END
END NOT
END LIBRARY

